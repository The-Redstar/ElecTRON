configuration countextend_behaviour_cfg of countextend is
   for behaviour
   end for;
end countextend_behaviour_cfg;
