configuration electron_synthesised_cfg of electron is
   for synthesised
   end for;
end electron_synthesised_cfg;
