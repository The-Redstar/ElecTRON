configuration pixelator_tb_behaviour_cfg of pixelator_tb is
   for behaviour
      for all: pixelator use configuration work.pixelator_behaviour_cfg;
      end for;
   end for;
end pixelator_tb_behaviour_cfg;
