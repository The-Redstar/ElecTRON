configuration memory_communication_behaviour_cfg of memory_communication is
   for behaviour
   end for;
end memory_communication_behaviour_cfg;
