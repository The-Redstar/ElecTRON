library IEEE;
use IEEE.std_logic_1164.ALL;

entity wall_decoder_tb is
end wall_decoder_tb;

