configuration memory_cntrll_behaviour_cfg of memory_cntrll is
   for behaviour
   end for;
end memory_cntrll_behaviour_cfg;
