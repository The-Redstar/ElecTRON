configuration engine_oscil_behaviour_cfg of engine_oscil is
   for behaviour
   end for;
end engine_oscil_behaviour_cfg;
