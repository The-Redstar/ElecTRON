configuration homescreen_behaviour_cfg of homescreen is
   for behaviour
   end for;
end homescreen_behaviour_cfg;
