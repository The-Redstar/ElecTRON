configuration flip_flop_behaviour_cfg of flip_flop is
   for behaviour
   end for;
end flip_flop_behaviour_cfg;
