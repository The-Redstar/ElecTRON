library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of ge_register_tb is
   component ge_register
   port(clk, reset	  : in  std_logic;	
   			e_position_0  : in  std_logic;
   			e_position_1  : in  std_logic;
   			d_position_0  : in  std_logic_vector(9 downto 0);
   			d_position_1  : in  std_logic_vector(9 downto 0);
   			e_layer_0	  : in  std_logic;		
   			e_layer_1	  : in  std_logic;
   			d_layer_0	  : in  std_logic;
   			d_layer_1	  : in  std_logic;
   			e_booster_0	  : in  std_logic;		
   			e_booster_1	  : in  std_logic;
   			d_booster_0	  : in  std_logic;
   			d_booster_1	  : in  std_logic;
   			e_boost_audio : in  std_logic;
   			d_boost_audio : in  std_logic_vector(1 downto 0);
   			e_booster_sync: in  std_logic;
   			d_booster_sync: in  std_logic;
   			e_next_layer_0: in  std_logic;
   			e_next_layer_1: in  std_logic;
   			d_next_layer_0: in  std_logic;
   			d_next_layer_1: in  std_logic;
   			e_border_0	  : in  std_logic;
   			e_border_1	  : in  std_logic;
   			d_border_0	  : in  std_logic;
   			d_border_1	  : in  std_logic;
   			e_read_mem    : in  std_logic;
   			d_read_mem    : in  std_logic_vector(7 downto 0);
   			e_direction_0 : in  std_logic;
   			e_direction_1 : in  std_logic;
   			d_direction_0 : in  std_logic_vector(1 downto 0);
   			d_direction_1 : in  std_logic_vector(1 downto 0);
   			e_next_dir_0  : in  std_logic;
   			e_next_dir_1  : in  std_logic;
   			d_next_dir_0  : in  std_logic_vector(1 downto 0);
   			d_next_dir_1  : in  std_logic_vector(1 downto 0);
   			e_p_state_0   : in  std_logic;
   			e_p_state_1   : in  std_logic;
   			d_p_state_0   : in  std_logic_vector(1 downto 0);
   			d_p_state_1   : in  std_logic_vector(1 downto 0);
   			e_map_select  : in  std_logic;
   			d_map_select  : in  std_logic_vector(1 downto 0);
   			e_speed_select: in  std_logic;
   			d_speed_select: in  std_logic_vector(1 downto 0);
   			q_position_0  : out std_logic_vector(9 downto 0);
   			q_position_1  : out std_logic_vector(9 downto 0);
   			q_layer_0	  : out std_logic;
   			q_layer_1	  : out std_logic;
   			q_booster_0	  : out std_logic;
   			q_booster_1	  : out std_logic;
   			q_boost_audio : out std_logic_vector(1 downto 0);
   			q_booster_sync	  : out std_logic;
   			q_next_layer_0: out std_logic;
   			q_next_layer_1: out std_logic;
   			q_border_0	  : out std_logic;
   			q_border_1	  : out std_logic;
   			q_read_mem    : out std_logic_vector(7 downto 0);
   			q_direction_0 : out std_logic_vector(1 downto 0);
   			q_direction_1 : out std_logic_vector(1 downto 0);
   			q_next_dir_0  : out std_logic_vector(1 downto 0);
   			q_next_dir_1  : out std_logic_vector(1 downto 0);
   			q_p_state_0   : out std_logic_vector(1 downto 0);
   			q_p_state_1   : out std_logic_vector(1 downto 0);
   			q_map_select  : out std_logic_vector(1 downto 0);
   			q_speed_select: out std_logic_vector(1 downto 0));
   end component;
   signal clk, reset	  : std_logic;
   signal e_position_0  : std_logic;
   signal e_position_1  : std_logic;
   signal d_position_0  : std_logic_vector(9 downto 0);
   signal d_position_1  : std_logic_vector(9 downto 0);
   signal e_layer_0	  : std_logic;
   signal e_layer_1	  : std_logic;
   signal d_layer_0	  : std_logic;
   signal d_layer_1	  : std_logic;
   signal e_booster_0	  : std_logic;
   signal e_booster_1	  : std_logic;
   signal d_booster_0	  : std_logic;
   signal d_booster_1	  : std_logic;
   signal e_boost_audio : std_logic;
   signal d_boost_audio : std_logic_vector(1 downto 0);
   signal e_booster_sync: std_logic;
   signal d_booster_sync: std_logic;
   signal e_next_layer_0: std_logic;
   signal e_next_layer_1: std_logic;
   signal d_next_layer_0: std_logic;
   signal d_next_layer_1: std_logic;
   signal e_border_0	  : std_logic;
   signal e_border_1	  : std_logic;
   signal d_border_0	  : std_logic;
   signal d_border_1	  : std_logic;
   signal e_read_mem    : std_logic;
   signal d_read_mem    : std_logic_vector(7 downto 0);
   signal e_direction_0 : std_logic;
   signal e_direction_1 : std_logic;
   signal d_direction_0 : std_logic_vector(1 downto 0);
   signal d_direction_1 : std_logic_vector(1 downto 0);
   signal e_next_dir_0  : std_logic;
   signal e_next_dir_1  : std_logic;
   signal d_next_dir_0  : std_logic_vector(1 downto 0);
   signal d_next_dir_1  : std_logic_vector(1 downto 0);
   signal e_p_state_0   : std_logic;
   signal e_p_state_1   : std_logic;
   signal d_p_state_0   : std_logic_vector(1 downto 0);
   signal d_p_state_1   : std_logic_vector(1 downto 0);
   signal e_map_select  : std_logic;
   signal d_map_select  : std_logic_vector(1 downto 0);
   signal e_speed_select: std_logic;
   signal d_speed_select: std_logic_vector(1 downto 0);
   signal q_position_0  : std_logic_vector(9 downto 0);
   signal q_position_1  : std_logic_vector(9 downto 0);
   signal q_layer_0	  : std_logic;
   signal q_layer_1	  : std_logic;
   signal q_booster_0	  : std_logic;
   signal q_booster_1	  : std_logic;
   signal q_boost_audio : std_logic_vector(1 downto 0);
   signal q_booster_sync	  : std_logic;
   signal q_next_layer_0: std_logic;
   signal q_next_layer_1: std_logic;
   signal q_border_0	  : std_logic;
   signal q_border_1	  : std_logic;
   signal q_read_mem    : std_logic_vector(7 downto 0);
   signal q_direction_0 : std_logic_vector(1 downto 0);
   signal q_direction_1 : std_logic_vector(1 downto 0);
   signal q_next_dir_0  : std_logic_vector(1 downto 0);
   signal q_next_dir_1  : std_logic_vector(1 downto 0);
   signal q_p_state_0   : std_logic_vector(1 downto 0);
   signal q_p_state_1   : std_logic_vector(1 downto 0);
   signal q_map_select  : std_logic_vector(1 downto 0);
   signal q_speed_select: std_logic_vector(1 downto 0);
begin
   test: ge_register port map (clk, reset, e_position_0, e_position_1, d_position_0, d_position_1, e_layer_0, e_layer_1, d_layer_0, d_layer_1, e_booster_0, e_booster_1, d_booster_0, d_booster_1, e_boost_audio, d_boost_audio, e_booster_sync, d_booster_sync, e_next_layer_0, e_next_layer_1, d_next_layer_0, d_next_layer_1, e_border_0, e_border_1, d_border_0, d_border_1, e_read_mem, d_read_mem, e_direction_0, e_direction_1, d_direction_0, d_direction_1, e_next_dir_0, e_next_dir_1, d_next_dir_0, d_next_dir_1, e_p_state_0, e_p_state_1, d_p_state_0, d_p_state_1, e_map_select, d_map_select, e_speed_select, d_speed_select, q_position_0, q_position_1, q_layer_0, q_layer_1, q_booster_0, q_booster_1, q_boost_audio, q_booster_sync, q_next_layer_0, q_next_layer_1, q_border_0, q_border_1, q_read_mem, q_direction_0, q_direction_1, q_next_dir_0, q_next_dir_1, q_p_state_0, q_p_state_1, q_map_select, q_speed_select);
   clk <= '0' after 0 ns,
          '1' after 20 ns when clk /= '1' else '0' after 20 ns;
   reset <= '1' after 0 ns,
            '0' after 80 ns;
   e_position_0 <= '0' after 0 ns, '1' after 100 ns, '0' after 140 ns;
   e_position_1 <= '0' after 0 ns, '1' after 200 ns, '0' after 240 ns;
   d_position_0(0) <= '1' after 0 ns;
   d_position_0(1) <= '0' after 0 ns;
   d_position_0(2) <= '0' after 0 ns;
   d_position_0(3) <= '0' after 0 ns;
   d_position_0(4) <= '0' after 0 ns;
   d_position_0(5) <= '0' after 0 ns;
   d_position_0(6) <= '0' after 0 ns;
   d_position_0(7) <= '0' after 0 ns;
   d_position_0(8) <= '0' after 0 ns;
   d_position_0(9) <= '0' after 0 ns;
   d_position_1(0) <= '1' after 0 ns;
   d_position_1(1) <= '0' after 0 ns;
   d_position_1(2) <= '0' after 0 ns;
   d_position_1(3) <= '0' after 0 ns;
   d_position_1(4) <= '0' after 0 ns;
   d_position_1(5) <= '0' after 0 ns;
   d_position_1(6) <= '0' after 0 ns;
   d_position_1(7) <= '0' after 0 ns;
   d_position_1(8) <= '0' after 0 ns;
   d_position_1(9) <= '0' after 0 ns;
   e_layer_0 <= '0' after 0 ns, '1' after 300 ns, '0' after 340 ns;
   e_layer_1 <= '0' after 0 ns, '1' after 400 ns, '0' after 440 ns;
   d_layer_0 <= '1' after 0 ns;
   d_layer_1 <= '1' after 0 ns;
   e_booster_0 <= '0' after 0 ns, '1' after 500 ns, '0' after 540 ns;
   e_booster_1 <= '0' after 0 ns, '1' after 600 ns, '0' after 640 ns;
   d_booster_0 <= '1' after 0 ns;
   d_booster_1 <= '1' after 0 ns;
   e_boost_audio <= '0' after 0 ns, '1' after 700 ns, '0' after 740 ns;
   d_boost_audio(0) <= '1' after 0 ns;
   d_boost_audio(1) <= '0' after 0 ns;
   e_booster_sync <= '0' after 0 ns, '1' after 800 ns, '0' after 840 ns;
   d_booster_sync <= '1' after 0 ns;
   e_next_layer_0 <= '0' after 0 ns, '1' after 900 ns, '0' after 940 ns;
   e_next_layer_1 <= '0' after 0 ns, '1' after 1000 ns, '0' after 1040 ns;
   d_next_layer_0 <= '1' after 0 ns;
   d_next_layer_1 <= '1' after 0 ns;
   e_border_0 <= '0' after 0 ns, '1' after 1100 ns, '0' after 1140 ns;
   e_border_1 <= '0' after 0 ns, '1' after 1200 ns, '0' after 1240 ns;
   d_border_0 <= '1' after 0 ns;
   d_border_1 <= '1' after 0 ns;
   e_read_mem <= '0' after 0 ns, '1' after 1300 ns, '0' after 1340 ns;
   d_read_mem(0) <= '1' after 0 ns;
   d_read_mem(1) <= '0' after 0 ns;
   d_read_mem(2) <= '0' after 0 ns;
   d_read_mem(3) <= '0' after 0 ns;
   d_read_mem(4) <= '0' after 0 ns;
   d_read_mem(5) <= '0' after 0 ns;
   d_read_mem(6) <= '0' after 0 ns;
   d_read_mem(7) <= '0' after 0 ns;
   e_direction_0 <= '0' after 0 ns, '1' after 1400 ns, '0' after 1440 ns;
   e_direction_1 <= '0' after 0 ns, '1' after 1500 ns, '0' after 1540 ns;
   d_direction_0(0) <= '1' after 0 ns;
   d_direction_0(1) <= '0' after 0 ns;
   d_direction_1(0) <= '1' after 0 ns;
   d_direction_1(1) <= '0' after 0 ns;
   e_next_dir_0 <= '0' after 0 ns, '1' after 1600 ns, '0' after 1640 ns;
   e_next_dir_1 <= '0' after 0 ns, '1' after 1700 ns, '0' after 1740 ns;
   d_next_dir_0(0) <= '1' after 0 ns;
   d_next_dir_0(1) <= '0' after 0 ns;
   d_next_dir_1(0) <= '1' after 0 ns;
   d_next_dir_1(1) <= '0' after 0 ns;
   e_p_state_0 <= '0' after 0 ns, '1' after 1800 ns, '0' after 1840 ns;
   e_p_state_1 <= '0' after 0 ns, '1' after 1900 ns, '0' after 1940 ns;
   d_p_state_0(0) <= '1' after 0 ns;
   d_p_state_0(1) <= '0' after 0 ns;
   d_p_state_1(0) <= '1' after 0 ns;
   d_p_state_1(1) <= '0' after 0 ns;
   e_map_select <= '0' after 0 ns, '1' after 2000 ns, '0' after 2040 ns;
   d_map_select(0) <= '1' after 0 ns;
   d_map_select(1) <= '0' after 0 ns;
   e_speed_select <= '0' after 0 ns, '1' after 2100 ns, '0' after 2140 ns;
   d_speed_select(0) <= '1' after 0 ns;
   d_speed_select(1) <= '0' after 0 ns;
end behaviour;

