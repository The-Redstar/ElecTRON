configuration color_bus_behaviour_cfg of color_bus is
   for behaviour
   end for;
end color_bus_behaviour_cfg;
