configuration pixelator_behaviour_cfg of pixelator is
   for behaviour
   end for;
end pixelator_behaviour_cfg;
