configuration memclear_behaviour_cfg of memclear is
   for behaviour
   end for;
end memclear_behaviour_cfg;
