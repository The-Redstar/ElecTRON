configuration wall_decoder_behaviour_cfg of wall_decoder is
   for behaviour
   end for;
end wall_decoder_behaviour_cfg;
