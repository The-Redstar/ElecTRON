configuration counter5b_tb_behaviour_cfg of counter5b_tb is
   for behaviour
      for all: counter5b use configuration work.counter5b_behaviour_cfg;
      end for;
   end for;
end counter5b_tb_behaviour_cfg;
