library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;

architecture behaviour of homescreen is

	signal x8_o100, y8_o56	: std_logic_vector(5 downto 0); --scaled down by a factor 8, offset
	signal x_o100,y_oc		: std_logic_vector(8 downto 0); --cycle offset to be finetuned
	signal y_o452,x_o208	: std_logic_vector(8 downto 0); --speed indicator offset
	
	
	type sprite_table is array (integer range <>,integer range <>) of std_logic;--index (y,x)
	
	constant logo_sprite1 : sprite_table(0 to 7, 0 to 63) := ("1111010000000000000000000000000000000000000000000000000000000000","1100010010001100000000000000000000000000000000000000000000000000","1110010111010000000000000000000000000000000000000000000000000000","1100010100010000000000000000000000000000000000000000000000000000","1111010010001100000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000");
	constant logo_sprite2 : sprite_table(0 to 7, 0 to 63) := ("0000000000000001111011100011001100100000000000000000000000000000","0000000000000000110011010110101110100000000000000000000000000000","0000000000000000110011100110101101100000000000000000000000000000","0000000000000000110011010110101100100000000000000000000000000000","0000000000000000110011010011001100100000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000");
	constant cycle_sprite : sprite_table(0 to 31, 0 to 255) := ("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000011111100000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000001110000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000011000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111110001111111111111111111111111000000000000001100000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111001100000001111111111111111000000000000000110000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111001100000000111111111111111000000000000000111000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000100000000111111111111111111111111111111111000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111100000100000000011111111111111111111001111111111000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111100000000011111111111111111100001111111111100000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111000111100000000011111111111111110000011110000111100000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110111100000001111111111111100000011000000001110000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111001110000010000001111111111111000000111000000001110000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001100000010000001111111111111000000110000000000110000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111001100000011111001111111111110000001110000000000110000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001100000000001111111111111110000001110000000000110000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111001100000000001111110000000001111111110000000000110000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110000000011110000000000000000000111000000001110000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111000110000000011100000000000000000000011000000001100000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111100001111000000000000000000000011110000111100000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111000000000000000000000011111111111100000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111000000000000000000000000000011111100000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000","0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
	constant speed_sprite_active : sprite_table(0 to 15, 0 to 15) := ("1111111110000000","0111111111000000","0011111111100000","0001111111110000","0000111111111000","0000011111111100","0000001111111110","0000000111111111","0000000111111111","0000001111111110","0000011111111100","0000111111111000","0001111111110000","0011111111100000","0111111111000000","1111111110000000");
	constant speed_sprite_inactive : sprite_table(0 to 15, 0 to 15) := ("1111111110000000","0110000011000000","0011000001100000","0001100000110000","0000110000011000","0000011000001100","0000001100000110","0000000110000011","0000000110000011","0000001100000110","0000011000001100","0000110000011000","0001100000110000","0011000001100000","0110000011000000","1111111110000000");

begin

	--coordinate signals
	x_o100	<= std_logic_vector(unsigned(x)-to_unsigned(100,9));
	x8_o100	<= x_o100(8 downto 3);
	y8_o56	<= std_logic_vector(unsigned(y(8 downto 3))-to_unsigned(7,6));
	y_oc	<= std_logic_vector(unsigned(y)-to_unsigned(110,9));
	y_o452	<= std_logic_vector(unsigned(y)-to_unsigned(452,9));
	x_o208	<= std_logic_vector(unsigned(x)-to_unsigned(208,9));



	process(x,y,pixelator,x_o100,x8_o100,y8_o56,y_oc)
		variable speed_pixel_active,speed_pixel_inactive: boolean;
	begin
		--default
		color <= "0000";
		
		--display logo
		--use scaled sprite, remove odd lines for effect
		if y(0)='0' and unsigned(y8_o56)<to_unsigned(8,5) then --and unsigned(x8_o56)<to_unsigned(8,5) then -> whitespace in sprite
			if logo_sprite1(to_integer(unsigned(y8_o56(2 downto 0))),to_integer(unsigned(x8_o100(5 downto 0))))='1' then
				color<="0011";
			elsif logo_sprite2(to_integer(unsigned(y8_o56(2 downto 0))),to_integer(unsigned(x8_o100(5 downto 0))))='1' then
				color<="1100";
			end if;
		end if;
		
		--display cycle
		if unsigned(y_oc)<to_unsigned(32,9) and x_o100(8)='0' then
			if cycle_sprite(to_integer(unsigned(y_oc(4 downto 0))),to_integer(unsigned(x_o100(7 downto 0))))='1' then
				color<="1111";
			end if;
		end if;
		
		--display scaled down map
		if to_unsigned(120,9)<=unsigned(x) and to_unsigned(200,9)<=unsigned(y) then
			if unsigned(x)<=to_unsigned(360,9) and unsigned(y)<=to_unsigned(440,9) then
				color<="1111";
			end if;
			if unsigned(x)<to_unsigned(360,9) and unsigned(y)<to_unsigned(440,9) then
				color<=pixelator;
			end if;
		end if;
		
		--display speed indicators
		speed_pixel_active	:=(  speed_sprite_active(to_integer(unsigned(y_o452(3 downto 0))),to_integer(unsigned(x_o208(3 downto 0))))='1');
		speed_pixel_inactive:=(speed_sprite_inactive(to_integer(unsigned(y_o452(3 downto 0))),to_integer(unsigned(x_o208(3 downto 0))))='1');
		if unsigned(y_o452)<to_unsigned(16,9) then
			if unsigned(x_o208)<to_unsigned(16,9) then
				if speed_pixel_active then
					color<="1111";
				end if;
			elsif unsigned(x_o208)<to_unsigned(32,9) then
				if speed_pixel_inactive or (speed_pixel_active and speed/="00") then
					color<="1111";
				end if;
			elsif unsigned(x_o208)<to_unsigned(48,9) then
				if speed_pixel_inactive or (speed_pixel_active and speed(1)='1') then
					color<="1111";
				end if;
			elsif unsigned(x_o208)<to_unsigned(64,9) then
				if speed_pixel_inactive or (speed_pixel_active and speed="11") then
					color<="1111";
				end if;
			end if;
		end if;
		
	end process;


end behaviour;

