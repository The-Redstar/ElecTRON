library IEEE;
use IEEE.std_logic_1164.ALL;

entity input_buffer_tb is
end input_buffer_tb;

