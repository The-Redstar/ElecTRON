configuration reg_10_behaviour_cfg of reg_10 is
   for behaviour
   end for;
end reg_10_behaviour_cfg;
