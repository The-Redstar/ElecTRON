library IEEE;
use IEEE.std_logic_1164.ALL;

entity memclear_tb is
end memclear_tb;

