configuration sidebar_tb_behaviour_cfg of sidebar_tb is
   for behaviour
      for all: sidebar use configuration work.sidebar_behaviour_cfg;
      end for;
   end for;
end sidebar_tb_behaviour_cfg;
