configuration readwrite_behaviour_cfg of readwrite is
   for behaviour
   end for;
end readwrite_behaviour_cfg;
