library IEEE;
use IEEE.std_logic_1164.ALL;

entity memory_cntrll_tb is
end memory_cntrll_tb;

