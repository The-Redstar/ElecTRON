configuration counter8b_behaviour_cfg of counter8b is
   for behaviour
   end for;
end counter8b_behaviour_cfg;
