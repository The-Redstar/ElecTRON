configuration counter8b_tb_behaviour_cfg of counter8b_tb is
   for behaviour
      for all: counter8b use configuration work.counter8b_behaviour_cfg;
      end for;
   end for;
end counter8b_tb_behaviour_cfg;
