library IEEE;
use IEEE.std_logic_1164.ALL;

entity grid_top_tb is
end grid_top_tb;

