library IEEE;
use IEEE.std_logic_1164.ALL;

entity pixelator_tb is
end pixelator_tb;

