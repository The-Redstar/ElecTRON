configuration electron_tb_behaviour_cfg of electron_tb is
   for behaviour
      for all: electron use configuration work.electron_structural_cfg;
      end for;
   end for;
end electron_tb_behaviour_cfg;
