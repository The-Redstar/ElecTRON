configuration memory_cntrll_tb_behaviour_cfg of memory_cntrll_tb is
   for behaviour
      for all: memory_cntrll use configuration work.memory_cntrll_behaviour_cfg;
      end for;
   end for;
end memory_cntrll_tb_behaviour_cfg;
