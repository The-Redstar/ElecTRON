
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture routed of electron is

  component DEL01BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL1BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD5BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD6BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component INVD2BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component XNR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKXOR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component MOAI22D1BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component CKAN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKXOR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component DFD0BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component DFKSND1BWP7T
    port(CP, D, SN : in std_logic; Q, QN : out std_logic);
  end component;

  component DFKSND0BWP7T
    port(CP, D, SN : in std_logic; Q, QN : out std_logic);
  end component;

  component IINR4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD5BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AO222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component OR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component AO32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component IIND4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component CKMUX2D1BWP7T
    port(I0, I1, S : in std_logic; Z : out std_logic);
  end component;

  component MUX2D1BWP7T
    port(I0, I1, S : in std_logic; Z : out std_logic);
  end component;

  component DFXQD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component HA1D0BWP7T
    port(A, B : in std_logic; CO, S : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component INR4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D1BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AO33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; Z : out std_logic);
  end component;

  component OAI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AN3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component OAI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OA31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component OA32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component OR4XD1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component AOI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component IND3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component OA32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AOI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component OA221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component OA22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component OA211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component OA33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; Z : out std_logic);
  end component;

  component AN2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OR3XD1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component AO31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component MAOI22D1BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AN3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component AOI21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AN4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component AN4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component MAOI222D1BWP7T
    port(A, B, C : in std_logic; ZN : out std_logic);
  end component;

  component MUX2ND0BWP7T
    port(I0, I1, S : in std_logic; ZN : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D1BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component FA1D0BWP7T
    port(A, B, CI : in std_logic; CO, S : out std_logic);
  end component;

  component NR3D1BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component EDFKCNQD1BWP7T
    port(CN, CP, D, E : in std_logic; Q : out std_logic);
  end component;

  component OR3D4BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component CKAN2D8BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OR4D4BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component DFCNQD1BWP7T
    port(CDN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component EDFCND1BWP7T
    port(CDN, CP, D, E : in std_logic; Q, QN : out std_logic);
  end component;

  component DFCND1BWP7T
    port(CDN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component OAI21D2BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OR3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  signal FE_PHN83_lbl1_rw_state_2, FE_PHN82_lbl0_mem_com_state_2, FE_PHN81_lbl0_border_0, FE_PHN80_lbl0_unsigned_busy_count_3, FE_PHN79_lbl1_rw_n_0 : std_logic;
  signal FE_PHN78_lbl0_n_62, FE_PHN77_lbl0_n_91, FE_PHN76_lbl1_rw_n_71, FE_PHN75_lbl0_n_110, FE_PHN74_lbl1_cex_n_6 : std_logic;
  signal FE_PHN73_lbl1_cey_n_6, FE_PHN72_lbl1_cm_n_24, FE_PHN71_lbl1_cey_n_3, FE_PHN70_lbl0_n_106, FE_PHN69_lbl1_rw_n_60 : std_logic;
  signal FE_PHN68_lbl1_cex_n_3, FE_PHN67_lbl0_n_107, FE_PHN66_lbl0_n_119, FE_PHN65_lbl0_n_117, FE_PHN64_read_memory_in_7 : std_logic;
  signal FE_PHN63_lbl2_v_count_9, FE_PHN62_lbl0_counter_busy_counter_state_1, FE_PHN61_lbl0_n_148, FE_PHN60_lbl0_booster_0, FE_PHN59_lbl0_next_layer_0 : std_logic;
  signal FE_PHN58_lbl0_next_direction_0_1, FE_PHN57_lbl0_unsigned_busy_count_6, FE_PHN56_lbl0_counter_busy_counter_state_0, FE_PHN55_lbl1_rw_n_29, FE_PHN54_lbl0_unsigned_busy_count_3 : std_logic;
  signal FE_PHN53_lbl1_ready_rw, FE_PHN52_lbl2_v_count_6, FE_PHN51_lbl0_border_0, FE_PHN50_lbl0_unsigned_busy_count_2, FE_PHN49_lbl0_unsigned_busy_count_1 : std_logic;
  signal FE_PHN48_lbl1_cm_n_23, FE_PHN47_lbl0_unsigned_busy_count_0, FE_PHN46_lbl0_booster_1, FE_PHN45_lbl2_v_count_7, FE_PHN44_lbl2_v_count_8 : std_logic;
  signal FE_PHN43_lbl1_cm_n_25, FE_PHN42_lbl0_border_1, FE_PHN41_lbl2_borders_synced_2, FE_PHN40_lbl1_cm_n_26, FE_PHN39_lbl0_next_direction_1_1 : std_logic;
  signal FE_PHN38_lbl2_data_synced_1, FE_PHN37_lbl1_cex_n_8, FE_PHN36_lbl0_mem_com_state_0, FE_PHN35_lbl2_borders_synced_7, FE_PHN34_read_memory_in_4 : std_logic;
  signal FE_PHN33_read_memory_in_5, FE_PHN32_read_memory_in_3, FE_PHN31_read_memory_in_2, FE_PHN30_lbl0_booster_sync, FE_PHN29_read_memory_in_0 : std_logic;
  signal FE_PHN28_read_memory_in_6, FE_PHN27_read_memory_in_1, FE_PHN26_lbl2_data_synced_5, FE_PHN25_lbl2_borders_synced_5, FE_PHN24_lbl2_jumps_synced_3 : std_logic;
  signal FE_PHN23_lbl2_data_synced_0, FE_PHN22_lbl2_jumps_synced_7, FE_PHN21_lbl2_data_synced_6, FE_PHN20_lbl2_borders_synced_6, FE_PHN19_lbl2_jumps_synced_5 : std_logic;
  signal FE_PHN18_lbl2_data_synced_2, FE_PHN17_lbl2_borders_synced_4, FE_PHN16_lbl2_jumps_synced_4, FE_PHN15_lbl2_jumps_synced_2, FE_PHN14_lbl2_borders_synced_3 : std_logic;
  signal FE_PHN13_lbl2_jumps_synced_0, FE_PHN12_lbl2_data_synced_4, FE_PHN11_lbl2_borders_synced_1, FE_PHN10_lbl2_borders_synced_0, FE_PHN9_lbl2_jumps_synced_6 : std_logic;
  signal FE_PHN8_lbl2_jumps_synced_1, FE_PHN7_lbl2_data_synced_7, FE_PHN6_lbl2_data_synced_3, FE_OFN5_memory_enable_out, FE_OFN4_lbl2_n_4 : std_logic;
  signal FE_OFN3_rst, CTS_12, CTS_11, FE_DBTN4_rst, FE_DBTN3_memory_reset_out : std_logic;
  signal FE_DBTN2_lbl2_h_count_3, FE_DBTN1_lbl2_h_count_1, FE_DBTN0_lbl2_v_count_2 : std_logic;
  signal position_1 : std_logic_vector(10 downto 0);
  signal position_0 : std_logic_vector(10 downto 0);
  signal lbl2_y_vec : std_logic_vector(4 downto 0);
  signal lbl2_central_x_vec : std_logic_vector(9 downto 0);
  signal lbl2_h_count : std_logic_vector(9 downto 0);
  signal lbl2_dx : std_logic_vector(3 downto 0);
  signal lbl2_v_count : std_logic_vector(9 downto 0);
  signal lbl2_dy_vec : std_logic_vector(3 downto 0);
  signal game_state : std_logic_vector(2 downto 0);
  signal lbl2_homescreen_color : std_logic_vector(3 downto 0);
  signal lbl2_pixelator_color : std_logic_vector(3 downto 0);
  signal lbl2_sidebar_color : std_logic_vector(3 downto 0);
  signal player_state_0 : std_logic_vector(1 downto 0);
  signal player_state_1 : std_logic_vector(1 downto 0);
  signal lbl2_borders_synced : std_logic_vector(7 downto 0);
  signal borders : std_logic_vector(7 downto 0);
  signal lbl2_data_synced : std_logic_vector(7 downto 0);
  signal lbl2_jumps_synced : std_logic_vector(7 downto 0);
  signal ramps : std_logic_vector(7 downto 0);
  signal lbl2_walls : std_logic_vector(7 downto 0);
  signal x_address : std_logic_vector(4 downto 0);
  signal start_position_0 : std_logic_vector(10 downto 0);
  signal y_address : std_logic_vector(4 downto 0);
  signal map_selected : std_logic_vector(1 downto 0);
  signal start_position_1 : std_logic_vector(10 downto 0);
  signal direction_1 : std_logic_vector(1 downto 0);
  signal direction_0 : std_logic_vector(1 downto 0);
  signal lbl0_d_position_1 : std_logic_vector(9 downto 0);
  signal address : std_logic_vector(9 downto 0);
  signal lbl0_next_direction_1 : std_logic_vector(1 downto 0);
  signal lbl0_next_direction_0 : std_logic_vector(1 downto 0);
  signal lbl0_d_position_0 : std_logic_vector(9 downto 0);
  signal lbl0_state : std_logic_vector(4 downto 0);
  signal write_memory : std_logic_vector(7 downto 0);
  signal lbl0_read_data_reg : std_logic_vector(7 downto 0);
  signal lbl0_d_read_data_reg : std_logic_vector(7 downto 0);
  signal lbl0_d_direction_0 : std_logic_vector(1 downto 0);
  signal lbl0_d_direction_1 : std_logic_vector(1 downto 0);
  signal lbl0_mem_com_state : std_logic_vector(3 downto 0);
  signal lbl0_d_next_direction_0 : std_logic_vector(1 downto 0);
  signal lbl0_d_next_direction_1 : std_logic_vector(1 downto 0);
  signal lbl0_d_speed_select : std_logic_vector(1 downto 0);
  signal lbl0_d_map_select : std_logic_vector(1 downto 0);
  signal lbl0_counter_busy_counter_state : std_logic_vector(1 downto 0);
  signal lbl0_unsigned_busy_count : std_logic_vector(6 downto 0);
  signal lbl1_cm_state : std_logic_vector(4 downto 0);
  signal lbl1_cex_state : std_logic_vector(1 downto 0);
  signal lbl1_rw_state : std_logic_vector(5 downto 0);
  signal lbl1_cur_w : std_logic_vector(7 downto 0);
  signal lbl1_cey_state : std_logic_vector(1 downto 0);
  signal UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2, UNCONNECTED3 : std_logic;
  signal UNCONNECTED4, busy, clear_memory, go_to, lbl0_booster_0 : std_logic;
  signal lbl0_booster_1, lbl0_booster_sync, lbl0_border_0, lbl0_border_1, lbl0_d_booster_0 : std_logic;
  signal lbl0_d_booster_1, lbl0_d_booster_sync, lbl0_d_layer_0, lbl0_d_layer_1, lbl0_e_position_0 : std_logic;
  signal lbl0_e_position_1, lbl0_mem_com_n_166, lbl0_mem_com_n_175, lbl0_n_0, lbl0_n_1 : std_logic;
  signal lbl0_n_4, lbl0_n_5, lbl0_n_6, lbl0_n_7, lbl0_n_8 : std_logic;
  signal lbl0_n_9, lbl0_n_10, lbl0_n_11, lbl0_n_12, lbl0_n_13 : std_logic;
  signal lbl0_n_14, lbl0_n_15, lbl0_n_16, lbl0_n_17, lbl0_n_18 : std_logic;
  signal lbl0_n_19, lbl0_n_20, lbl0_n_21, lbl0_n_22, lbl0_n_23 : std_logic;
  signal lbl0_n_25, lbl0_n_26, lbl0_n_27, lbl0_n_28, lbl0_n_29 : std_logic;
  signal lbl0_n_30, lbl0_n_31, lbl0_n_32, lbl0_n_33, lbl0_n_34 : std_logic;
  signal lbl0_n_35, lbl0_n_36, lbl0_n_37, lbl0_n_38, lbl0_n_39 : std_logic;
  signal lbl0_n_40, lbl0_n_41, lbl0_n_43, lbl0_n_44, lbl0_n_45 : std_logic;
  signal lbl0_n_46, lbl0_n_47, lbl0_n_48, lbl0_n_49, lbl0_n_50 : std_logic;
  signal lbl0_n_51, lbl0_n_52, lbl0_n_53, lbl0_n_54, lbl0_n_55 : std_logic;
  signal lbl0_n_56, lbl0_n_57, lbl0_n_58, lbl0_n_60, lbl0_n_61 : std_logic;
  signal lbl0_n_62, lbl0_n_63, lbl0_n_64, lbl0_n_65, lbl0_n_66 : std_logic;
  signal lbl0_n_67, lbl0_n_68, lbl0_n_69, lbl0_n_70, lbl0_n_71 : std_logic;
  signal lbl0_n_72, lbl0_n_73, lbl0_n_74, lbl0_n_75, lbl0_n_76 : std_logic;
  signal lbl0_n_77, lbl0_n_78, lbl0_n_79, lbl0_n_80, lbl0_n_81 : std_logic;
  signal lbl0_n_82, lbl0_n_83, lbl0_n_84, lbl0_n_85, lbl0_n_86 : std_logic;
  signal lbl0_n_87, lbl0_n_88, lbl0_n_89, lbl0_n_90, lbl0_n_91 : std_logic;
  signal lbl0_n_92, lbl0_n_93, lbl0_n_94, lbl0_n_95, lbl0_n_96 : std_logic;
  signal lbl0_n_97, lbl0_n_98, lbl0_n_99, lbl0_n_100, lbl0_n_101 : std_logic;
  signal lbl0_n_102, lbl0_n_103, lbl0_n_104, lbl0_n_105, lbl0_n_106 : std_logic;
  signal lbl0_n_107, lbl0_n_108, lbl0_n_109, lbl0_n_110, lbl0_n_111 : std_logic;
  signal lbl0_n_112, lbl0_n_113, lbl0_n_114, lbl0_n_115, lbl0_n_116 : std_logic;
  signal lbl0_n_117, lbl0_n_118, lbl0_n_119, lbl0_n_120, lbl0_n_121 : std_logic;
  signal lbl0_n_122, lbl0_n_123, lbl0_n_124, lbl0_n_125, lbl0_n_126 : std_logic;
  signal lbl0_n_127, lbl0_n_128, lbl0_n_129, lbl0_n_130, lbl0_n_131 : std_logic;
  signal lbl0_n_132, lbl0_n_133, lbl0_n_134, lbl0_n_135, lbl0_n_136 : std_logic;
  signal lbl0_n_137, lbl0_n_138, lbl0_n_139, lbl0_n_140, lbl0_n_141 : std_logic;
  signal lbl0_n_142, lbl0_n_143, lbl0_n_144, lbl0_n_145, lbl0_n_147 : std_logic;
  signal lbl0_n_148, lbl0_n_149, lbl0_n_150, lbl0_n_151, lbl0_n_152 : std_logic;
  signal lbl0_n_153, lbl0_n_154, lbl0_n_155, lbl0_n_156, lbl0_n_157 : std_logic;
  signal lbl0_n_158, lbl0_n_159, lbl0_n_160, lbl0_n_161, lbl0_n_162 : std_logic;
  signal lbl0_n_163, lbl0_n_164, lbl0_n_165, lbl0_n_166, lbl0_n_167 : std_logic;
  signal lbl0_n_168, lbl0_n_169, lbl0_n_170, lbl0_n_171, lbl0_n_172 : std_logic;
  signal lbl0_n_173, lbl0_n_174, lbl0_n_175, lbl0_n_176, lbl0_n_177 : std_logic;
  signal lbl0_n_178, lbl0_n_179, lbl0_n_180, lbl0_n_181, lbl0_n_182 : std_logic;
  signal lbl0_n_183, lbl0_n_184, lbl0_n_185, lbl0_n_186, lbl0_n_187 : std_logic;
  signal lbl0_n_188, lbl0_n_189, lbl0_n_190, lbl0_n_191, lbl0_n_192 : std_logic;
  signal lbl0_n_193, lbl0_n_194, lbl0_n_195, lbl0_n_196, lbl0_n_197 : std_logic;
  signal lbl0_n_198, lbl0_n_199, lbl0_n_200, lbl0_n_201, lbl0_n_202 : std_logic;
  signal lbl0_n_203, lbl0_n_204, lbl0_n_205, lbl0_n_206, lbl0_n_207 : std_logic;
  signal lbl0_n_208, lbl0_n_209, lbl0_n_210, lbl0_n_211, lbl0_n_212 : std_logic;
  signal lbl0_n_213, lbl0_n_214, lbl0_n_215, lbl0_n_216, lbl0_n_217 : std_logic;
  signal lbl0_n_218, lbl0_n_219, lbl0_n_220, lbl0_n_221, lbl0_n_222 : std_logic;
  signal lbl0_n_223, lbl0_n_224, lbl0_n_225, lbl0_n_226, lbl0_n_227 : std_logic;
  signal lbl0_n_228, lbl0_n_229, lbl0_n_230, lbl0_n_231, lbl0_n_232 : std_logic;
  signal lbl0_n_233, lbl0_n_234, lbl0_n_235, lbl0_n_236, lbl0_n_237 : std_logic;
  signal lbl0_n_238, lbl0_n_239, lbl0_n_240, lbl0_n_241, lbl0_n_242 : std_logic;
  signal lbl0_n_243, lbl0_n_244, lbl0_n_245, lbl0_n_246, lbl0_n_247 : std_logic;
  signal lbl0_n_248, lbl0_n_249, lbl0_n_250, lbl0_n_251, lbl0_n_252 : std_logic;
  signal lbl0_n_253, lbl0_n_254, lbl0_n_255, lbl0_n_256, lbl0_n_257 : std_logic;
  signal lbl0_n_258, lbl0_n_259, lbl0_n_260, lbl0_n_261, lbl0_n_262 : std_logic;
  signal lbl0_n_263, lbl0_n_264, lbl0_n_265, lbl0_n_266, lbl0_n_267 : std_logic;
  signal lbl0_n_268, lbl0_n_269, lbl0_n_270, lbl0_n_271, lbl0_n_272 : std_logic;
  signal lbl0_n_273, lbl0_n_274, lbl0_n_275, lbl0_n_276, lbl0_n_277 : std_logic;
  signal lbl0_n_278, lbl0_n_279, lbl0_n_280, lbl0_n_281, lbl0_n_282 : std_logic;
  signal lbl0_n_283, lbl0_n_284, lbl0_n_285, lbl0_n_286, lbl0_n_287 : std_logic;
  signal lbl0_n_288, lbl0_n_289, lbl0_n_290, lbl0_n_291, lbl0_n_292 : std_logic;
  signal lbl0_n_293, lbl0_n_294, lbl0_n_295, lbl0_n_296, lbl0_n_297 : std_logic;
  signal lbl0_n_298, lbl0_n_299, lbl0_n_300, lbl0_n_301, lbl0_n_302 : std_logic;
  signal lbl0_n_303, lbl0_n_304, lbl0_n_305, lbl0_n_306, lbl0_n_307 : std_logic;
  signal lbl0_n_308, lbl0_n_309, lbl0_n_310, lbl0_n_311, lbl0_n_312 : std_logic;
  signal lbl0_n_313, lbl0_n_314, lbl0_n_315, lbl0_n_316, lbl0_n_317 : std_logic;
  signal lbl0_n_318, lbl0_n_319, lbl0_n_320, lbl0_n_321, lbl0_n_322 : std_logic;
  signal lbl0_n_323, lbl0_n_324, lbl0_n_325, lbl0_n_326, lbl0_n_327 : std_logic;
  signal lbl0_n_328, lbl0_n_329, lbl0_n_330, lbl0_n_331, lbl0_n_332 : std_logic;
  signal lbl0_n_333, lbl0_n_334, lbl0_n_335, lbl0_n_336, lbl0_n_337 : std_logic;
  signal lbl0_n_338, lbl0_n_339, lbl0_n_340, lbl0_n_341, lbl0_n_342 : std_logic;
  signal lbl0_n_343, lbl0_n_344, lbl0_n_345, lbl0_n_346, lbl0_n_347 : std_logic;
  signal lbl0_n_348, lbl0_n_349, lbl0_n_350, lbl0_n_351, lbl0_n_352 : std_logic;
  signal lbl0_n_353, lbl0_n_354, lbl0_n_355, lbl0_n_356, lbl0_n_357 : std_logic;
  signal lbl0_n_358, lbl0_n_359, lbl0_n_360, lbl0_n_361, lbl0_n_362 : std_logic;
  signal lbl0_n_363, lbl0_n_364, lbl0_n_365, lbl0_n_366, lbl0_n_367 : std_logic;
  signal lbl0_n_368, lbl0_n_369, lbl0_n_370, lbl0_n_371, lbl0_n_372 : std_logic;
  signal lbl0_n_373, lbl0_n_374, lbl0_n_375, lbl0_n_376, lbl0_n_377 : std_logic;
  signal lbl0_n_378, lbl0_n_379, lbl0_n_380, lbl0_n_381, lbl0_n_382 : std_logic;
  signal lbl0_n_383, lbl0_n_384, lbl0_n_385, lbl0_n_386, lbl0_n_387 : std_logic;
  signal lbl0_n_388, lbl0_n_389, lbl0_n_390, lbl0_n_391, lbl0_n_392 : std_logic;
  signal lbl0_n_393, lbl0_n_394, lbl0_n_395, lbl0_n_396, lbl0_n_397 : std_logic;
  signal lbl0_n_398, lbl0_n_399, lbl0_n_400, lbl0_n_401, lbl0_n_402 : std_logic;
  signal lbl0_n_403, lbl0_n_404, lbl0_n_405, lbl0_n_406, lbl0_n_407 : std_logic;
  signal lbl0_n_408, lbl0_n_410, lbl0_n_411, lbl0_n_412, lbl0_n_413 : std_logic;
  signal lbl0_n_414, lbl0_n_415, lbl0_n_416, lbl0_n_417, lbl0_n_418 : std_logic;
  signal lbl0_n_419, lbl0_n_420, lbl0_n_421, lbl0_n_422, lbl0_n_423 : std_logic;
  signal lbl0_n_424, lbl0_n_425, lbl0_n_426, lbl0_n_427, lbl0_n_428 : std_logic;
  signal lbl0_n_429, lbl0_n_430, lbl0_n_432, lbl0_n_433, lbl0_n_436 : std_logic;
  signal lbl0_n_437, lbl0_n_471, lbl0_n_472, lbl0_n_473, lbl0_n_474 : std_logic;
  signal lbl0_n_476, lbl0_n_477, lbl0_n_504, lbl0_n_505, lbl0_n_506 : std_logic;
  signal lbl0_n_507, lbl0_n_508, lbl0_n_509, lbl0_n_510, lbl0_n_511 : std_logic;
  signal lbl0_n_512, lbl0_n_513, lbl0_n_515, lbl0_n_516, lbl0_n_517 : std_logic;
  signal lbl0_n_1952_BAR, lbl0_next_layer_0, lbl0_next_layer_1, lbl1_cex_n_2, lbl1_cex_n_3 : std_logic;
  signal lbl1_cex_n_4, lbl1_cex_n_5, lbl1_cex_n_6, lbl1_cex_n_7, lbl1_cex_n_8 : std_logic;
  signal lbl1_cex_n_9, lbl1_cey_n_2, lbl1_cey_n_3, lbl1_cey_n_4, lbl1_cey_n_5 : std_logic;
  signal lbl1_cey_n_6, lbl1_cey_n_7, lbl1_cey_n_8, lbl1_cey_n_9, lbl1_clr_rst : std_logic;
  signal lbl1_cm_n_2, lbl1_cm_n_3, lbl1_cm_n_4, lbl1_cm_n_5, lbl1_cm_n_6 : std_logic;
  signal lbl1_cm_n_7, lbl1_cm_n_8, lbl1_cm_n_9, lbl1_cm_n_10, lbl1_cm_n_11 : std_logic;
  signal lbl1_cm_n_12, lbl1_cm_n_13, lbl1_cm_n_14, lbl1_cm_n_15, lbl1_cm_n_16 : std_logic;
  signal lbl1_cm_n_17, lbl1_cm_n_18, lbl1_cm_n_20, lbl1_cm_n_21, lbl1_cm_n_22 : std_logic;
  signal lbl1_cm_n_23, lbl1_cm_n_24, lbl1_cm_n_25, lbl1_cm_n_26, lbl1_cm_n_27 : std_logic;
  signal lbl1_cm_n_28, lbl1_cm_n_29, lbl1_cm_n_32, lbl1_cm_n_37, lbl1_cm_n_52 : std_logic;
  signal lbl1_cw_n_0, lbl1_cw_n_2, lbl1_cw_n_3, lbl1_cw_n_4, lbl1_cw_n_5 : std_logic;
  signal lbl1_cw_n_6, lbl1_cw_n_7, lbl1_cw_n_8, lbl1_cw_n_9, lbl1_cw_n_10 : std_logic;
  signal lbl1_cw_n_11, lbl1_cw_n_12, lbl1_cw_n_13, lbl1_cw_n_14, lbl1_cx_n_0 : std_logic;
  signal lbl1_cx_n_2, lbl1_cx_n_3, lbl1_cx_n_4, lbl1_cx_n_5, lbl1_cx_n_6 : std_logic;
  signal lbl1_cx_n_7, lbl1_cx_n_8, lbl1_cy_n_0, lbl1_cy_n_2, lbl1_cy_n_3 : std_logic;
  signal lbl1_cy_n_4, lbl1_cy_n_5, lbl1_cy_n_6, lbl1_cy_n_7, lbl1_cy_n_8 : std_logic;
  signal lbl1_me_clr, lbl1_me_rw, lbl1_n_1, lbl1_ready_clr, lbl1_ready_rw : std_logic;
  signal lbl1_rw_n_0, lbl1_rw_n_3, lbl1_rw_n_4, lbl1_rw_n_5, lbl1_rw_n_6 : std_logic;
  signal lbl1_rw_n_7, lbl1_rw_n_8, lbl1_rw_n_9, lbl1_rw_n_10, lbl1_rw_n_11 : std_logic;
  signal lbl1_rw_n_12, lbl1_rw_n_13, lbl1_rw_n_14, lbl1_rw_n_15, lbl1_rw_n_16 : std_logic;
  signal lbl1_rw_n_17, lbl1_rw_n_18, lbl1_rw_n_19, lbl1_rw_n_20, lbl1_rw_n_21 : std_logic;
  signal lbl1_rw_n_22, lbl1_rw_n_23, lbl1_rw_n_24, lbl1_rw_n_25, lbl1_rw_n_26 : std_logic;
  signal lbl1_rw_n_27, lbl1_rw_n_28, lbl1_rw_n_29, lbl1_rw_n_30, lbl1_rw_n_31 : std_logic;
  signal lbl1_rw_n_32, lbl1_rw_n_33, lbl1_rw_n_34, lbl1_rw_n_35, lbl1_rw_n_36 : std_logic;
  signal lbl1_rw_n_37, lbl1_rw_n_38, lbl1_rw_n_39, lbl1_rw_n_40, lbl1_rw_n_41 : std_logic;
  signal lbl1_rw_n_42, lbl1_rw_n_43, lbl1_rw_n_44, lbl1_rw_n_45, lbl1_rw_n_46 : std_logic;
  signal lbl1_rw_n_47, lbl1_rw_n_48, lbl1_rw_n_49, lbl1_rw_n_50, lbl1_rw_n_51 : std_logic;
  signal lbl1_rw_n_52, lbl1_rw_n_53, lbl1_rw_n_54, lbl1_rw_n_55, lbl1_rw_n_56 : std_logic;
  signal lbl1_rw_n_57, lbl1_rw_n_58, lbl1_rw_n_59, lbl1_rw_n_60, lbl1_rw_n_61 : std_logic;
  signal lbl1_rw_n_62, lbl1_rw_n_63, lbl1_rw_n_64, lbl1_rw_n_65, lbl1_rw_n_66 : std_logic;
  signal lbl1_rw_n_67, lbl1_rw_n_68, lbl1_rw_n_69, lbl1_rw_n_70, lbl1_rw_n_71 : std_logic;
  signal lbl1_rw_n_72, lbl1_rw_n_73, lbl1_rw_n_74, lbl1_rw_n_75, lbl1_rw_n_76 : std_logic;
  signal lbl1_rw_n_77, lbl1_rw_n_78, lbl1_rw_n_79, lbl1_rw_n_80, lbl1_rw_n_81 : std_logic;
  signal lbl1_rw_n_82, lbl1_rw_n_83, lbl1_rw_n_84, lbl1_rw_n_85, lbl1_rw_n_86 : std_logic;
  signal lbl1_rw_n_87, lbl1_rw_n_88, lbl1_rw_n_89, lbl1_rw_n_90, lbl1_rw_n_97 : std_logic;
  signal lbl1_rw_n_99, lbl1_rw_n_100, lbl1_rw_rst, lbl1_we_clr, lbl1_we_rw : std_logic;
  signal lbl1_x_incr1, lbl1_x_incr2, lbl1_x_incr3, lbl1_y_incr1, lbl1_y_incr2 : std_logic;
  signal lbl1_y_incr3, lbl2_dec0_n_0, lbl2_dec0_n_1, lbl2_dec0_n_2, lbl2_dec0_n_3 : std_logic;
  signal lbl2_dec0_n_5, lbl2_dec1_n_0, lbl2_dec1_n_1, lbl2_dec1_n_2, lbl2_dec1_n_3 : std_logic;
  signal lbl2_dec1_n_5, lbl2_hscr_n_0, lbl2_hscr_n_1, lbl2_hscr_n_2, lbl2_hscr_n_3 : std_logic;
  signal lbl2_hscr_n_6, lbl2_hscr_n_9, lbl2_hscr_n_10, lbl2_hscr_n_11, lbl2_hscr_n_12 : std_logic;
  signal lbl2_hscr_n_13, lbl2_hscr_n_14, lbl2_hscr_n_15, lbl2_hscr_n_16, lbl2_hscr_n_17 : std_logic;
  signal lbl2_hscr_n_18, lbl2_hscr_n_19, lbl2_hscr_n_20, lbl2_hscr_n_21, lbl2_hscr_n_22 : std_logic;
  signal lbl2_hscr_n_23, lbl2_hscr_n_24, lbl2_hscr_n_25, lbl2_hscr_n_26, lbl2_hscr_n_27 : std_logic;
  signal lbl2_hscr_n_28, lbl2_hscr_n_29, lbl2_hscr_n_30, lbl2_hscr_n_31, lbl2_hscr_n_32 : std_logic;
  signal lbl2_hscr_n_33, lbl2_hscr_n_34, lbl2_hscr_n_35, lbl2_hscr_n_36, lbl2_hscr_n_37 : std_logic;
  signal lbl2_hscr_n_38, lbl2_hscr_n_39, lbl2_hscr_n_40, lbl2_hscr_n_41, lbl2_hscr_n_42 : std_logic;
  signal lbl2_hscr_n_43, lbl2_hscr_n_44, lbl2_hscr_n_45, lbl2_hscr_n_46, lbl2_hscr_n_47 : std_logic;
  signal lbl2_hscr_n_48, lbl2_hscr_n_49, lbl2_hscr_n_50, lbl2_hscr_n_51, lbl2_hscr_n_52 : std_logic;
  signal lbl2_hscr_n_53, lbl2_hscr_n_54, lbl2_hscr_n_55, lbl2_hscr_n_56, lbl2_hscr_n_57 : std_logic;
  signal lbl2_hscr_n_58, lbl2_hscr_n_59, lbl2_hscr_n_60, lbl2_hscr_n_61, lbl2_hscr_n_62 : std_logic;
  signal lbl2_hscr_n_63, lbl2_hscr_n_64, lbl2_hscr_n_65, lbl2_hscr_n_66, lbl2_hscr_n_67 : std_logic;
  signal lbl2_hscr_n_68, lbl2_hscr_n_70, lbl2_hscr_n_71, lbl2_hscr_n_72, lbl2_hscr_n_73 : std_logic;
  signal lbl2_hscr_n_74, lbl2_hscr_n_76, lbl2_hscr_n_77, lbl2_hscr_n_78, lbl2_hscr_n_79 : std_logic;
  signal lbl2_hscr_n_80, lbl2_hscr_n_81, lbl2_hscr_n_82, lbl2_hscr_n_83, lbl2_hscr_n_84 : std_logic;
  signal lbl2_hscr_n_85, lbl2_hscr_n_86, lbl2_hscr_n_87, lbl2_hscr_n_88, lbl2_hscr_n_89 : std_logic;
  signal lbl2_hscr_n_90, lbl2_hscr_n_91, lbl2_hscr_n_92, lbl2_hscr_n_93, lbl2_hscr_n_94 : std_logic;
  signal lbl2_hscr_n_95, lbl2_hscr_n_96, lbl2_hscr_n_97, lbl2_hscr_n_98, lbl2_hscr_n_99 : std_logic;
  signal lbl2_hscr_n_100, lbl2_hscr_n_101, lbl2_hscr_n_102, lbl2_hscr_n_103, lbl2_hscr_n_104 : std_logic;
  signal lbl2_hscr_n_105, lbl2_hscr_n_106, lbl2_hscr_n_107, lbl2_hscr_n_108, lbl2_hscr_n_109 : std_logic;
  signal lbl2_hscr_n_110, lbl2_hscr_n_111, lbl2_hscr_n_112, lbl2_hscr_n_113, lbl2_hscr_n_114 : std_logic;
  signal lbl2_hscr_n_115, lbl2_hscr_n_116, lbl2_hscr_n_117, lbl2_hscr_n_118, lbl2_hscr_n_119 : std_logic;
  signal lbl2_hscr_n_120, lbl2_hscr_n_121, lbl2_hscr_n_122, lbl2_hscr_n_123, lbl2_hscr_n_124 : std_logic;
  signal lbl2_hscr_n_125, lbl2_hscr_n_126, lbl2_hscr_n_127, lbl2_hscr_n_128, lbl2_hscr_n_129 : std_logic;
  signal lbl2_hscr_n_130, lbl2_hscr_n_131, lbl2_hscr_n_132, lbl2_hscr_n_133, lbl2_hscr_n_134 : std_logic;
  signal lbl2_hscr_n_135, lbl2_hscr_n_136, lbl2_hscr_n_137, lbl2_hscr_n_138, lbl2_hscr_n_139 : std_logic;
  signal lbl2_hscr_n_140, lbl2_hscr_n_141, lbl2_hscr_n_142, lbl2_hscr_n_143, lbl2_hscr_n_144 : std_logic;
  signal lbl2_hscr_n_145, lbl2_hscr_n_146, lbl2_hscr_n_147, lbl2_hscr_n_148, lbl2_hscr_n_149 : std_logic;
  signal lbl2_hscr_n_150, lbl2_hscr_n_151, lbl2_hscr_n_153, lbl2_hscr_n_154, lbl2_hscr_n_155 : std_logic;
  signal lbl2_hscr_n_156, lbl2_hscr_n_157, lbl2_hscr_n_158, lbl2_hscr_n_159, lbl2_hscr_n_160 : std_logic;
  signal lbl2_hscr_n_161, lbl2_hscr_n_162, lbl2_hscr_n_163, lbl2_hscr_n_164, lbl2_hscr_n_165 : std_logic;
  signal lbl2_hscr_n_166, lbl2_hscr_n_167, lbl2_hscr_n_168, lbl2_hscr_n_169, lbl2_hscr_n_170 : std_logic;
  signal lbl2_hscr_n_171, lbl2_hscr_n_172, lbl2_hscr_n_173, lbl2_hscr_n_174, lbl2_hscr_n_175 : std_logic;
  signal lbl2_hscr_n_176, lbl2_hscr_n_177, lbl2_hscr_n_178, lbl2_hscr_n_179, lbl2_hscr_n_180 : std_logic;
  signal lbl2_hscr_n_181, lbl2_hscr_n_182, lbl2_hscr_n_183, lbl2_hscr_n_184, lbl2_hscr_n_185 : std_logic;
  signal lbl2_hscr_n_186, lbl2_hscr_n_187, lbl2_hscr_n_188, lbl2_hscr_n_189, lbl2_hscr_n_190 : std_logic;
  signal lbl2_hscr_n_191, lbl2_hscr_n_192, lbl2_hscr_n_193, lbl2_hscr_n_194, lbl2_hscr_n_195 : std_logic;
  signal lbl2_hscr_n_196, lbl2_hscr_n_197, lbl2_hscr_n_198, lbl2_hscr_n_199, lbl2_hscr_n_200 : std_logic;
  signal lbl2_hscr_n_201, lbl2_hscr_n_202, lbl2_hscr_n_203, lbl2_hscr_n_204, lbl2_hscr_n_205 : std_logic;
  signal lbl2_hscr_n_206, lbl2_hscr_n_207, lbl2_hscr_n_208, lbl2_hscr_n_209, lbl2_hscr_n_210 : std_logic;
  signal lbl2_hscr_n_211, lbl2_hscr_n_212, lbl2_hscr_n_213, lbl2_hscr_n_214, lbl2_hscr_n_215 : std_logic;
  signal lbl2_hscr_n_216, lbl2_hscr_n_217, lbl2_hscr_n_218, lbl2_hscr_n_219, lbl2_hscr_n_220 : std_logic;
  signal lbl2_hscr_n_221, lbl2_hscr_n_222, lbl2_hscr_n_223, lbl2_hscr_n_224, lbl2_hscr_n_225 : std_logic;
  signal lbl2_hscr_n_226, lbl2_hscr_n_227, lbl2_hscr_n_228, lbl2_hscr_n_229, lbl2_hscr_n_230 : std_logic;
  signal lbl2_hscr_n_231, lbl2_hscr_n_232, lbl2_hscr_n_233, lbl2_hscr_n_234, lbl2_hscr_n_235 : std_logic;
  signal lbl2_hscr_n_236, lbl2_hscr_n_237, lbl2_hscr_n_238, lbl2_hscr_n_239, lbl2_hscr_n_240 : std_logic;
  signal lbl2_hscr_n_241, lbl2_hscr_n_242, lbl2_hscr_n_243, lbl2_hscr_n_244, lbl2_hscr_n_245 : std_logic;
  signal lbl2_hscr_n_246, lbl2_hscr_n_247, lbl2_hscr_n_248, lbl2_hscr_n_249, lbl2_hscr_n_250 : std_logic;
  signal lbl2_hscr_n_251, lbl2_hscr_n_252, lbl2_hscr_n_253, lbl2_hscr_n_254, lbl2_hscr_n_255 : std_logic;
  signal lbl2_hscr_n_256, lbl2_hscr_n_257, lbl2_hscr_n_258, lbl2_hscr_n_259, lbl2_hscr_n_260 : std_logic;
  signal lbl2_hscr_n_261, lbl2_hscr_n_262, lbl2_hscr_n_263, lbl2_hscr_n_264, lbl2_hscr_n_265 : std_logic;
  signal lbl2_hscr_n_266, lbl2_hscr_n_267, lbl2_hscr_n_268, lbl2_hscr_n_269, lbl2_hscr_n_270 : std_logic;
  signal lbl2_hscr_n_271, lbl2_hscr_n_272, lbl2_hscr_n_273, lbl2_hscr_n_274, lbl2_hscr_n_275 : std_logic;
  signal lbl2_hscr_n_276, lbl2_hscr_n_277, lbl2_hscr_n_278, lbl2_hscr_n_279, lbl2_hscr_n_280 : std_logic;
  signal lbl2_hscr_n_281, lbl2_hscr_n_282, lbl2_hscr_n_283, lbl2_hscr_n_284, lbl2_hscr_n_285 : std_logic;
  signal lbl2_hscr_n_286, lbl2_hscr_n_287, lbl2_hscr_n_288, lbl2_hscr_n_289, lbl2_hscr_n_290 : std_logic;
  signal lbl2_hscr_n_291, lbl2_hscr_n_292, lbl2_hscr_n_293, lbl2_hscr_n_294, lbl2_hscr_n_295 : std_logic;
  signal lbl2_hscr_n_296, lbl2_hscr_n_297, lbl2_hscr_n_298, lbl2_hscr_n_299, lbl2_hscr_n_300 : std_logic;
  signal lbl2_hscr_n_301, lbl2_hscr_n_302, lbl2_hscr_n_303, lbl2_hscr_n_304, lbl2_hscr_n_305 : std_logic;
  signal lbl2_hscr_n_306, lbl2_hscr_n_307, lbl2_hscr_n_308, lbl2_hscr_n_309, lbl2_hscr_n_310 : std_logic;
  signal lbl2_hscr_n_311, lbl2_hscr_n_312, lbl2_hscr_n_313, lbl2_hscr_n_314, lbl2_hscr_n_315 : std_logic;
  signal lbl2_hscr_n_316, lbl2_hscr_n_317, lbl2_hscr_n_318, lbl2_hscr_n_319, lbl2_hscr_n_320 : std_logic;
  signal lbl2_hscr_n_321, lbl2_hscr_n_322, lbl2_hscr_n_323, lbl2_hscr_n_324, lbl2_hscr_n_325 : std_logic;
  signal lbl2_hscr_n_326, lbl2_hscr_n_327, lbl2_hscr_n_328, lbl2_hscr_n_329, lbl2_hscr_n_330 : std_logic;
  signal lbl2_hscr_n_331, lbl2_hscr_n_332, lbl2_hscr_n_333, lbl2_hscr_n_334, lbl2_hscr_n_335 : std_logic;
  signal lbl2_hscr_n_336, lbl2_hscr_n_337, lbl2_hscr_n_338, lbl2_hscr_n_339, lbl2_hscr_n_340 : std_logic;
  signal lbl2_hscr_n_341, lbl2_hscr_n_342, lbl2_hscr_n_343, lbl2_hscr_n_344, lbl2_hscr_n_345 : std_logic;
  signal lbl2_hscr_n_346, lbl2_hscr_n_347, lbl2_hscr_n_348, lbl2_hscr_n_349, lbl2_hscr_n_350 : std_logic;
  signal lbl2_hscr_n_351, lbl2_hscr_n_352, lbl2_hscr_n_353, lbl2_hscr_n_354, lbl2_hscr_n_355 : std_logic;
  signal lbl2_hscr_n_356, lbl2_hscr_n_357, lbl2_hscr_n_358, lbl2_hscr_n_359, lbl2_hscr_n_360 : std_logic;
  signal lbl2_hscr_n_361, lbl2_hscr_n_362, lbl2_hscr_n_363, lbl2_hscr_n_364, lbl2_hscr_n_365 : std_logic;
  signal lbl2_hscr_n_366, lbl2_hscr_n_367, lbl2_hscr_n_368, lbl2_hscr_n_369, lbl2_hscr_n_370 : std_logic;
  signal lbl2_hscr_n_371, lbl2_hscr_n_400, lbl2_hscr_n_401, lbl2_n_2, lbl2_n_3 : std_logic;
  signal lbl2_n_4, lbl2_n_5, lbl2_n_6, lbl2_n_7, lbl2_n_8 : std_logic;
  signal lbl2_n_9, lbl2_n_10, lbl2_n_11, lbl2_n_12, lbl2_n_13 : std_logic;
  signal lbl2_n_14, lbl2_n_15, lbl2_n_16, lbl2_n_17, lbl2_n_18 : std_logic;
  signal lbl2_n_19, lbl2_n_20, lbl2_n_21, lbl2_n_22, lbl2_n_23 : std_logic;
  signal lbl2_n_24, lbl2_n_25, lbl2_n_26, lbl2_n_27, lbl2_n_28 : std_logic;
  signal lbl2_n_29, lbl2_n_30, lbl2_n_31, lbl2_n_32, lbl2_n_33 : std_logic;
  signal lbl2_n_34, lbl2_n_35, lbl2_n_36, lbl2_n_37, lbl2_n_38 : std_logic;
  signal lbl2_n_39, lbl2_n_40, lbl2_n_41, lbl2_n_42, lbl2_n_43 : std_logic;
  signal lbl2_n_44, lbl2_n_45, lbl2_n_46, lbl2_n_47, lbl2_n_48 : std_logic;
  signal lbl2_n_49, lbl2_n_50, lbl2_n_51, lbl2_n_52, lbl2_n_53 : std_logic;
  signal lbl2_n_56, lbl2_n_58, lbl2_n_59, lbl2_n_65, lbl2_n_66 : std_logic;
  signal lbl2_n_67, lbl2_n_68, lbl2_n_69, lbl2_n_70, lbl2_n_71 : std_logic;
  signal lbl2_n_72, lbl2_n_73, lbl2_n_74, lbl2_n_75, lbl2_n_76 : std_logic;
  signal lbl2_n_78, lbl2_n_79, lbl2_n_80, lbl2_n_82, lbl2_n_83 : std_logic;
  signal lbl2_n_84, lbl2_n_85, lbl2_n_86, lbl2_n_87, lbl2_n_88 : std_logic;
  signal lbl2_n_89, lbl2_n_90, lbl2_n_91, lbl2_n_92, lbl2_n_93 : std_logic;
  signal lbl2_n_94, lbl2_n_95, lbl2_n_96, lbl2_n_97, lbl2_n_98 : std_logic;
  signal lbl2_n_99, lbl2_n_100, lbl2_n_101, lbl2_n_102, lbl2_n_103 : std_logic;
  signal lbl2_n_104, lbl2_n_105, lbl2_n_106, lbl2_n_107, lbl2_n_108 : std_logic;
  signal lbl2_n_109, lbl2_n_110, lbl2_n_111, lbl2_n_112, lbl2_n_114 : std_logic;
  signal lbl2_n_115, lbl2_n_116, lbl2_n_117, lbl2_n_118, lbl2_n_119 : std_logic;
  signal lbl2_n_120, lbl2_n_121, lbl2_n_123, lbl2_n_124, lbl2_n_125 : std_logic;
  signal lbl2_n_126, lbl2_n_127, lbl2_n_128, lbl2_n_129, lbl2_n_130 : std_logic;
  signal lbl2_n_131, lbl2_n_132, lbl2_n_133, lbl2_n_134, lbl2_n_135 : std_logic;
  signal lbl2_n_136, lbl2_n_137, lbl2_n_138, lbl2_n_139, lbl2_n_140 : std_logic;
  signal lbl2_n_141, lbl2_n_142, lbl2_n_143, lbl2_n_146, lbl2_n_147 : std_logic;
  signal lbl2_n_148, lbl2_n_149, lbl2_n_150, lbl2_n_151, lbl2_n_152 : std_logic;
  signal lbl2_n_153, lbl2_n_154, lbl2_n_156, lbl2_n_158, lbl2_n_189 : std_logic;
  signal lbl2_n_190, lbl2_n_225, lbl2_n_226, lbl2_n_227, lbl2_pxl_n_0 : std_logic;
  signal lbl2_pxl_n_1, lbl2_pxl_n_2, lbl2_pxl_n_3, lbl2_pxl_n_4, lbl2_pxl_n_5 : std_logic;
  signal lbl2_pxl_n_6, lbl2_pxl_n_7, lbl2_pxl_n_8, lbl2_pxl_n_9, lbl2_pxl_n_10 : std_logic;
  signal lbl2_pxl_n_11, lbl2_pxl_n_12, lbl2_pxl_n_13, lbl2_pxl_n_14, lbl2_pxl_n_15 : std_logic;
  signal lbl2_pxl_n_16, lbl2_pxl_n_17, lbl2_pxl_n_18, lbl2_pxl_n_19, lbl2_pxl_n_20 : std_logic;
  signal lbl2_pxl_n_21, lbl2_pxl_n_22, lbl2_pxl_n_23, lbl2_pxl_n_24, lbl2_pxl_n_25 : std_logic;
  signal lbl2_pxl_n_26, lbl2_pxl_n_27, lbl2_pxl_n_28, lbl2_pxl_n_29, lbl2_pxl_n_30 : std_logic;
  signal lbl2_pxl_n_31, lbl2_pxl_n_32, lbl2_pxl_n_33, lbl2_pxl_n_34, lbl2_pxl_n_35 : std_logic;
  signal lbl2_pxl_n_36, lbl2_pxl_n_37, lbl2_pxl_n_38, lbl2_pxl_n_39, lbl2_pxl_n_40 : std_logic;
  signal lbl2_pxl_n_41, lbl2_pxl_n_42, lbl2_pxl_n_43, lbl2_pxl_n_44, lbl2_pxl_n_45 : std_logic;
  signal lbl2_pxl_n_46, lbl2_pxl_n_47, lbl2_pxl_n_48, lbl2_pxl_n_49, lbl2_pxl_n_50 : std_logic;
  signal lbl2_pxl_n_51, lbl2_pxl_n_52, lbl2_pxl_n_53, lbl2_pxl_n_54, lbl2_pxl_n_55 : std_logic;
  signal lbl2_pxl_n_56, lbl2_pxl_n_57, lbl2_pxl_n_58, lbl2_pxl_n_59, lbl2_pxl_n_60 : std_logic;
  signal lbl2_pxl_n_61, lbl2_pxl_n_62, lbl2_pxl_n_63, lbl2_pxl_n_64, lbl2_pxl_n_65 : std_logic;
  signal lbl2_pxl_n_66, lbl2_pxl_n_67, lbl2_pxl_n_68, lbl2_pxl_n_69, lbl2_pxl_n_70 : std_logic;
  signal lbl2_pxl_n_71, lbl2_pxl_n_72, lbl2_pxl_n_73, lbl2_pxl_n_74, lbl2_pxl_n_75 : std_logic;
  signal lbl2_pxl_n_76, lbl2_pxl_n_77, lbl2_pxl_n_78, lbl2_pxl_n_79, lbl2_pxl_n_80 : std_logic;
  signal lbl2_pxl_n_81, lbl2_pxl_n_82, lbl2_pxl_n_83, lbl2_pxl_n_84, lbl2_pxl_n_85 : std_logic;
  signal lbl2_pxl_n_86, lbl2_pxl_n_87, lbl2_pxl_n_88, lbl2_pxl_n_89, lbl2_pxl_n_90 : std_logic;
  signal lbl2_pxl_n_91, lbl2_pxl_n_92, lbl2_pxl_n_93, lbl2_pxl_n_94, lbl2_pxl_n_95 : std_logic;
  signal lbl2_pxl_n_96, lbl2_pxl_n_97, lbl2_pxl_n_98, lbl2_pxl_n_99, lbl2_pxl_n_100 : std_logic;
  signal lbl2_pxl_n_101, lbl2_pxl_n_102, lbl2_pxl_n_103, lbl2_pxl_n_104, lbl2_pxl_n_105 : std_logic;
  signal lbl2_pxl_n_106, lbl2_pxl_n_107, lbl2_pxl_n_108, lbl2_pxl_n_109, lbl2_pxl_n_110 : std_logic;
  signal lbl2_pxl_n_111, lbl2_pxl_n_112, lbl2_pxl_n_113, lbl2_pxl_n_114, lbl2_pxl_n_115 : std_logic;
  signal lbl2_pxl_n_116, lbl2_pxl_n_117, lbl2_pxl_n_118, lbl2_pxl_n_119, lbl2_pxl_n_120 : std_logic;
  signal lbl2_pxl_n_121, lbl2_pxl_n_122, lbl2_pxl_n_123, lbl2_pxl_n_124, lbl2_pxl_n_125 : std_logic;
  signal lbl2_pxl_n_126, lbl2_pxl_n_127, lbl2_pxl_n_128, lbl2_pxl_n_129, lbl2_pxl_n_130 : std_logic;
  signal lbl2_pxl_n_131, lbl2_pxl_n_132, lbl2_pxl_n_133, lbl2_pxl_n_134, lbl2_pxl_n_135 : std_logic;
  signal lbl2_pxl_n_136, lbl2_pxl_n_137, lbl2_pxl_n_138, lbl2_pxl_n_139, lbl2_pxl_n_140 : std_logic;
  signal lbl2_pxl_n_141, lbl2_pxl_n_142, lbl2_pxl_n_143, lbl2_pxl_n_144, lbl2_pxl_n_145 : std_logic;
  signal lbl2_pxl_n_146, lbl2_pxl_n_147, lbl2_pxl_n_148, lbl2_pxl_n_149, lbl2_pxl_n_150 : std_logic;
  signal lbl2_pxl_n_151, lbl2_pxl_n_152, lbl2_pxl_n_153, lbl2_pxl_n_154, lbl2_pxl_n_155 : std_logic;
  signal lbl2_pxl_n_156, lbl2_pxl_n_157, lbl2_pxl_n_158, lbl2_pxl_n_159, lbl2_pxl_n_160 : std_logic;
  signal lbl2_pxl_n_161, lbl2_pxl_n_162, lbl2_pxl_n_163, lbl2_pxl_n_164, lbl2_pxl_n_165 : std_logic;
  signal lbl2_pxl_n_166, lbl2_pxl_n_167, lbl2_pxl_n_168, lbl2_pxl_n_169, lbl2_pxl_n_170 : std_logic;
  signal lbl2_pxl_n_171, lbl2_pxl_n_172, lbl2_pxl_n_173, lbl2_pxl_n_174, lbl2_pxl_n_175 : std_logic;
  signal lbl2_pxl_n_176, lbl2_pxl_n_177, lbl2_pxl_n_178, lbl2_pxl_n_179, lbl2_pxl_n_180 : std_logic;
  signal lbl2_pxl_n_181, lbl2_pxl_n_182, lbl2_pxl_n_183, lbl2_pxl_n_184, lbl2_pxl_n_185 : std_logic;
  signal lbl2_pxl_n_186, lbl2_pxl_n_187, lbl2_pxl_n_188, lbl2_pxl_n_189, lbl2_pxl_n_190 : std_logic;
  signal lbl2_pxl_n_191, lbl2_pxl_n_192, lbl2_pxl_n_193, lbl2_pxl_n_194, lbl2_pxl_n_195 : std_logic;
  signal lbl2_pxl_n_196, lbl2_pxl_n_197, lbl2_pxl_n_198, lbl2_pxl_n_199, lbl2_pxl_n_200 : std_logic;
  signal lbl2_pxl_n_201, lbl2_pxl_n_202, lbl2_pxl_n_203, lbl2_pxl_n_205, lbl2_pxl_n_206 : std_logic;
  signal lbl2_pxl_n_207, lbl2_pxl_n_208, lbl2_pxl_n_210, lbl2_sdb_n_0, lbl2_sdb_n_2 : std_logic;
  signal lbl2_sdb_n_5, lbl2_sdb_n_6, lbl2_sdb_n_7, lbl2_sdb_n_8, lbl2_sdb_n_9 : std_logic;
  signal lbl2_sdb_n_10, lbl2_sdb_n_11, lbl2_sdb_n_12, lbl2_sdb_n_13, lbl2_sdb_n_14 : std_logic;
  signal lbl2_sdb_n_15, lbl2_sdb_n_16, lbl2_sdb_n_17, lbl2_sdb_n_18, lbl2_sdb_n_19 : std_logic;
  signal lbl2_sdb_n_20, lbl2_sdb_n_21, lbl2_sdb_n_22, lbl2_sdb_n_23, lbl2_sdb_n_24 : std_logic;
  signal lbl2_sdb_n_25, lbl2_sdb_n_26, lbl2_sdb_n_27, lbl2_sdb_n_28, lbl2_sdb_n_29 : std_logic;
  signal lbl2_sdb_n_30, lbl2_sdb_n_31, lbl2_sdb_n_32, lbl2_sdb_n_33, lbl2_sdb_n_34 : std_logic;
  signal lbl2_sdb_n_35, lbl2_sdb_n_36, lbl2_sdb_n_37, lbl2_sdb_n_38, lbl2_sdb_n_39 : std_logic;
  signal lbl2_sdb_n_40, lbl2_sdb_n_41, lbl2_sdb_n_42, lbl2_sdb_n_43, lbl2_sdb_n_44 : std_logic;
  signal lbl2_sdb_n_45, lbl2_sdb_n_46, lbl2_sdb_n_47, lbl2_sdb_n_48, lbl2_sdb_n_49 : std_logic;
  signal lbl2_sdb_n_50, lbl2_sdb_n_51, lbl2_sdb_n_52, lbl2_sdb_n_53, lbl2_sdb_n_54 : std_logic;
  signal lbl2_sdb_n_55, lbl2_sdb_n_56, lbl2_sdb_n_57, lbl2_sdb_n_58, lbl2_sdb_n_59 : std_logic;
  signal lbl2_sdb_n_60, lbl2_sdb_n_61, lbl2_sdb_n_62, lbl2_sdb_n_63, lbl2_sdb_n_64 : std_logic;
  signal lbl2_sdb_n_65, lbl2_sdb_n_66, lbl2_sdb_n_67, lbl2_sdb_n_68, lbl2_sdb_n_69 : std_logic;
  signal lbl2_sdb_n_70, lbl2_sdb_n_71, lbl2_sdb_n_72, lbl2_sdb_n_73, lbl2_sdb_n_74 : std_logic;
  signal lbl2_sdb_n_75, lbl2_sdb_n_76, lbl2_sdb_n_77, lbl2_sdb_n_78, lbl2_sdb_n_79 : std_logic;
  signal lbl2_sdb_n_80, lbl2_sdb_n_81, lbl2_sdb_n_82, lbl2_sdb_n_83, lbl2_sdb_n_84 : std_logic;
  signal lbl2_sdb_n_85, lbl2_sdb_n_86, lbl2_sdb_n_87, lbl2_sdb_n_88, lbl2_sdb_n_89 : std_logic;
  signal lbl2_sdb_n_90, lbl2_sdb_n_91, lbl2_sdb_n_92, lbl2_sdb_n_93, lbl2_sdb_n_94 : std_logic;
  signal lbl2_sdb_n_95, lbl2_sdb_n_96, lbl2_sdb_n_97, lbl2_sdb_n_98, lbl2_sdb_n_99 : std_logic;
  signal lbl2_sdb_n_100, lbl2_sdb_n_101, lbl2_sdb_n_102, lbl2_sdb_n_103, lbl2_sdb_n_104 : std_logic;
  signal lbl2_sdb_n_105, lbl2_sdb_n_106, lbl2_sdb_n_107, lbl2_sdb_n_108, lbl2_sdb_n_109 : std_logic;
  signal lbl2_sdb_n_110, lbl2_sdb_n_111, lbl2_sdb_n_112, lbl2_sdb_n_113, lbl2_sdb_n_114 : std_logic;
  signal lbl2_sdb_n_115, lbl2_sdb_n_116, lbl2_sdb_n_117, lbl2_sdb_n_118, lbl2_sdb_n_119 : std_logic;
  signal lbl2_sdb_n_120, lbl2_sdb_n_121, lbl2_sdb_n_122, lbl2_sdb_n_123, lbl2_sdb_n_124 : std_logic;
  signal lbl2_sdb_n_125, lbl2_sdb_n_126, lbl2_sdb_n_127, lbl2_sdb_n_128, lbl2_sdb_n_129 : std_logic;
  signal lbl2_sdb_n_130, lbl2_sdb_n_131, lbl2_sdb_n_132, lbl2_sdb_n_133, lbl2_sdb_n_134 : std_logic;
  signal lbl2_sdb_n_135, lbl2_sdb_n_136, lbl2_sdb_n_137, lbl2_sdb_n_138, lbl2_sdb_n_139 : std_logic;
  signal lbl2_sdb_n_140, lbl2_sdb_n_141, lbl2_sdb_n_142, lbl2_sdb_n_143, lbl2_sdb_n_144 : std_logic;
  signal lbl2_sdb_n_145, lbl2_sdb_n_146, lbl2_sdb_n_147, lbl2_sdb_n_148, lbl2_sdb_n_149 : std_logic;
  signal lbl2_sdb_n_150, lbl2_sdb_n_151, lbl2_sdb_n_152, lbl2_sdb_n_153, lbl2_sdb_n_154 : std_logic;
  signal lbl2_sdb_n_155, lbl2_sdb_n_156, lbl2_sdb_n_157, lbl2_sdb_n_158, lbl2_sdb_n_159 : std_logic;
  signal lbl2_sdb_n_160, lbl2_sdb_n_161, lbl2_sdb_n_162, lbl2_sdb_n_163, lbl2_sdb_n_164 : std_logic;
  signal lbl2_sdb_n_165, lbl2_sdb_n_166, lbl2_sdb_n_167, lbl2_sdb_n_168, lbl2_sdb_n_169 : std_logic;
  signal lbl2_sdb_n_170, lbl2_sdb_n_171, lbl2_sdb_n_172, lbl2_sdb_n_173, lbl2_sdb_n_174 : std_logic;
  signal lbl2_sdb_n_175, lbl2_sdb_n_176, lbl2_sdb_n_177, lbl2_sdb_n_178, lbl2_sdb_n_179 : std_logic;
  signal lbl4_n_3, lbl4_n_4, lbl4_n_5, lbl4_n_6, lbl4_n_7 : std_logic;
  signal lbl4_n_8, lbl4_n_9, lbl4_n_11, lbl4_n_12, lbl4_n_13 : std_logic;
  signal lbl4_n_14, lbl4_n_15, lbl4_n_16, lbl4_n_17, lbl4_n_18 : std_logic;
  signal lbl4_n_19, lbl4_n_20, lbl4_n_21, lbl4_n_22, lbl4_n_23 : std_logic;
  signal lbl4_n_25, lbl4_n_26, lbl4_n_27, lbl4_n_29, lbl4_n_30 : std_logic;
  signal lbl4_n_31, lbl4_n_32, lbl4_n_33, lbl4_n_34, lbl4_n_35 : std_logic;
  signal lbl4_n_36, lbl4_n_37, lbl4_n_38, lbl4_n_40, lbl4_n_41 : std_logic;
  signal lbl4_n_42, lbl4_n_43, lbl4_n_44, lbl4_n_45, lbl4_n_46 : std_logic;
  signal lbl4_n_47, lbl4_n_48, lbl4_n_49, lbl4_n_50, lbl4_n_51 : std_logic;
  signal lbl4_n_52, lbl4_n_53, lbl4_n_54, lbl4_n_55, lbl4_n_56 : std_logic;
  signal lbl4_n_57, lbl4_n_58, lbl4_n_59, lbl4_n_60, lbl4_n_61 : std_logic;
  signal lbl4_n_62, lbl4_n_63, lbl4_n_64, lbl4_n_65, lbl4_n_66 : std_logic;
  signal lbl4_n_67, lbl4_n_68, lbl4_n_69, lbl4_n_70, lbl4_n_71 : std_logic;
  signal lbl4_n_72, lbl4_n_73, lbl4_n_74, lbl4_n_75, lbl4_n_76 : std_logic;
  signal lbl4_n_77, lbl4_n_78, lbl4_n_79, lbl4_n_80, lbl4_n_81 : std_logic;
  signal lbl4_n_82, lbl4_n_83, lbl4_n_84, lbl4_n_86, lbl4_n_87 : std_logic;
  signal lbl4_n_88, lbl4_n_89, lbl4_n_90, lbl4_n_91, lbl4_n_92 : std_logic;
  signal lbl4_n_93, lbl4_n_94, lbl4_n_95, lbl4_n_96, lbl4_n_97 : std_logic;
  signal lbl4_n_98, lbl4_n_99, lbl4_n_100, lbl4_n_101, lbl4_n_102 : std_logic;
  signal lbl4_n_103, lbl4_n_104, lbl4_n_105, lbl4_n_106, lbl4_n_107 : std_logic;
  signal lbl4_n_108, lbl4_n_109, lbl4_n_110, lbl4_n_111, lbl4_n_112 : std_logic;
  signal lbl4_n_113, lbl4_n_114, lbl4_n_115, lbl4_n_116, lbl4_n_117 : std_logic;
  signal lbl4_n_118, lbl4_n_121, lbl4_n_122, lbl4_n_123, lbl4_n_124 : std_logic;
  signal lbl4_n_125, lbl4_n_126, lbl4_n_127, lbl4_n_129, lbl4_n_131 : std_logic;
  signal lbl4_n_132, lbl4_n_134, lbl4_n_138, lbl4_n_139, lbl4_n_142 : std_logic;
  signal lbl4_n_161, memory_ready, reset_vga_mem, write_enable, x_increment : std_logic;
  signal y_increment : std_logic;

begin

  FE_PHC83_lbl1_rw_state_2 : DEL01BWP7T port map(I => lbl1_rw_state(2), Z => FE_PHN83_lbl1_rw_state_2);
  FE_PHC82_lbl0_mem_com_state_2 : DEL01BWP7T port map(I => lbl0_mem_com_state(2), Z => FE_PHN82_lbl0_mem_com_state_2);
  FE_PHC81_lbl0_border_0 : DEL01BWP7T port map(I => lbl0_border_0, Z => FE_PHN81_lbl0_border_0);
  FE_PHC80_lbl0_unsigned_busy_count_3 : BUFFD3BWP7T port map(I => lbl0_unsigned_busy_count(3), Z => FE_PHN80_lbl0_unsigned_busy_count_3);
  FE_PHC79_lbl1_rw_n_0 : CKBD0BWP7T port map(I => lbl1_rw_n_0, Z => FE_PHN79_lbl1_rw_n_0);
  FE_PHC78_lbl0_n_62 : CKBD0BWP7T port map(I => FE_PHN78_lbl0_n_62, Z => lbl0_n_62);
  FE_PHC77_lbl0_n_91 : DEL01BWP7T port map(I => lbl0_n_91, Z => FE_PHN77_lbl0_n_91);
  FE_PHC76_lbl1_rw_n_71 : DEL0BWP7T port map(I => lbl1_rw_n_71, Z => FE_PHN76_lbl1_rw_n_71);
  FE_PHC75_lbl0_n_110 : DEL0BWP7T port map(I => FE_PHN75_lbl0_n_110, Z => lbl0_n_110);
  FE_PHC74_lbl1_cex_n_6 : DEL0BWP7T port map(I => lbl1_cex_n_6, Z => FE_PHN74_lbl1_cex_n_6);
  FE_PHC73_lbl1_cey_n_6 : DEL0BWP7T port map(I => lbl1_cey_n_6, Z => FE_PHN73_lbl1_cey_n_6);
  FE_PHC72_lbl1_cm_n_24 : DEL0BWP7T port map(I => lbl1_cm_n_24, Z => FE_PHN72_lbl1_cm_n_24);
  FE_PHC71_lbl1_cey_n_3 : DEL1BWP7T port map(I => FE_PHN71_lbl1_cey_n_3, Z => lbl1_cey_n_3);
  FE_PHC70_lbl0_n_106 : DEL2BWP7T port map(I => lbl0_n_106, Z => FE_PHN70_lbl0_n_106);
  FE_PHC69_lbl1_rw_n_60 : DEL0BWP7T port map(I => lbl1_rw_n_60, Z => FE_PHN69_lbl1_rw_n_60);
  FE_PHC68_lbl1_cex_n_3 : DEL0BWP7T port map(I => lbl1_cex_n_3, Z => FE_PHN68_lbl1_cex_n_3);
  FE_PHC67_lbl0_n_107 : DEL1BWP7T port map(I => lbl0_n_107, Z => FE_PHN67_lbl0_n_107);
  FE_PHC66_lbl0_n_119 : DEL1BWP7T port map(I => FE_PHN66_lbl0_n_119, Z => lbl0_n_119);
  FE_PHC65_lbl0_n_117 : DEL1BWP7T port map(I => lbl0_n_117, Z => FE_PHN65_lbl0_n_117);
  FE_PHC64_read_memory_in_7 : DEL0BWP7T port map(I => read_memory_in(7), Z => FE_PHN64_read_memory_in_7);
  FE_PHC63_lbl2_v_count_9 : DEL0BWP7T port map(I => FE_PHN63_lbl2_v_count_9, Z => lbl2_v_count(9));
  FE_PHC62_lbl0_counter_busy_counter_state_1 : DEL0BWP7T port map(I => FE_PHN62_lbl0_counter_busy_counter_state_1, Z => lbl0_counter_busy_counter_state(1));
  FE_PHC61_lbl0_n_148 : DEL01BWP7T port map(I => lbl0_n_148, Z => FE_PHN61_lbl0_n_148);
  FE_PHC60_lbl0_booster_0 : DEL0BWP7T port map(I => lbl0_booster_0, Z => FE_PHN60_lbl0_booster_0);
  FE_PHC59_lbl0_next_layer_0 : DEL01BWP7T port map(I => lbl0_next_layer_0, Z => FE_PHN59_lbl0_next_layer_0);
  FE_PHC58_lbl0_next_direction_0_1 : DEL01BWP7T port map(I => lbl0_next_direction_0(1), Z => FE_PHN58_lbl0_next_direction_0_1);
  FE_PHC57_lbl0_unsigned_busy_count_6 : DEL1BWP7T port map(I => FE_PHN57_lbl0_unsigned_busy_count_6, Z => lbl0_unsigned_busy_count(6));
  FE_PHC56_lbl0_counter_busy_counter_state_0 : DEL1BWP7T port map(I => FE_PHN56_lbl0_counter_busy_counter_state_0, Z => lbl0_counter_busy_counter_state(0));
  FE_PHC55_lbl1_rw_n_29 : BUFFD3BWP7T port map(I => lbl1_rw_n_29, Z => FE_PHN55_lbl1_rw_n_29);
  FE_PHC54_lbl0_unsigned_busy_count_3 : DEL0BWP7T port map(I => FE_PHN54_lbl0_unsigned_busy_count_3, Z => lbl0_unsigned_busy_count(3));
  FE_PHC53_lbl1_ready_rw : DEL0BWP7T port map(I => lbl1_ready_rw, Z => FE_PHN53_lbl1_ready_rw);
  FE_PHC52_lbl2_v_count_6 : CKBD0BWP7T port map(I => lbl2_v_count(6), Z => FE_PHN52_lbl2_v_count_6);
  FE_PHC51_lbl0_border_0 : CKBD0BWP7T port map(I => FE_PHN81_lbl0_border_0, Z => FE_PHN51_lbl0_border_0);
  FE_PHC50_lbl0_unsigned_busy_count_2 : DEL1BWP7T port map(I => lbl0_unsigned_busy_count(2), Z => FE_PHN50_lbl0_unsigned_busy_count_2);
  FE_PHC49_lbl0_unsigned_busy_count_1 : DEL1BWP7T port map(I => FE_PHN49_lbl0_unsigned_busy_count_1, Z => lbl0_unsigned_busy_count(1));
  FE_PHC48_lbl1_cm_n_23 : DEL0BWP7T port map(I => FE_PHN48_lbl1_cm_n_23, Z => lbl1_cm_n_23);
  FE_PHC47_lbl0_unsigned_busy_count_0 : DEL1BWP7T port map(I => FE_PHN47_lbl0_unsigned_busy_count_0, Z => lbl0_unsigned_busy_count(0));
  FE_PHC46_lbl0_booster_1 : DEL01BWP7T port map(I => lbl0_booster_1, Z => FE_PHN46_lbl0_booster_1);
  FE_PHC45_lbl2_v_count_7 : CKBD0BWP7T port map(I => lbl2_v_count(7), Z => FE_PHN45_lbl2_v_count_7);
  FE_PHC44_lbl2_v_count_8 : CKBD0BWP7T port map(I => lbl2_v_count(8), Z => FE_PHN44_lbl2_v_count_8);
  FE_PHC43_lbl1_cm_n_25 : DEL0BWP7T port map(I => lbl1_cm_n_25, Z => FE_PHN43_lbl1_cm_n_25);
  FE_PHC42_lbl0_border_1 : DEL0BWP7T port map(I => lbl0_border_1, Z => FE_PHN42_lbl0_border_1);
  FE_PHC41_lbl2_borders_synced_2 : DEL1BWP7T port map(I => lbl2_borders_synced(2), Z => FE_PHN41_lbl2_borders_synced_2);
  FE_PHC40_lbl1_cm_n_26 : DEL0BWP7T port map(I => lbl1_cm_n_26, Z => FE_PHN40_lbl1_cm_n_26);
  FE_PHC39_lbl0_next_direction_1_1 : CKBD0BWP7T port map(I => lbl0_next_direction_1(1), Z => FE_PHN39_lbl0_next_direction_1_1);
  FE_PHC38_lbl2_data_synced_1 : DEL1BWP7T port map(I => lbl2_data_synced(1), Z => FE_PHN38_lbl2_data_synced_1);
  FE_PHC37_lbl1_cex_n_8 : DEL0BWP7T port map(I => lbl1_cex_n_8, Z => FE_PHN37_lbl1_cex_n_8);
  FE_PHC36_lbl0_mem_com_state_0 : DEL0BWP7T port map(I => lbl0_mem_com_state(0), Z => FE_PHN36_lbl0_mem_com_state_0);
  FE_PHC35_lbl2_borders_synced_7 : DEL2BWP7T port map(I => lbl2_borders_synced(7), Z => FE_PHN35_lbl2_borders_synced_7);
  FE_PHC34_read_memory_in_4 : CKBD0BWP7T port map(I => read_memory_in(4), Z => FE_PHN34_read_memory_in_4);
  FE_PHC33_read_memory_in_5 : CKBD0BWP7T port map(I => read_memory_in(5), Z => FE_PHN33_read_memory_in_5);
  FE_PHC32_read_memory_in_3 : CKBD0BWP7T port map(I => read_memory_in(3), Z => FE_PHN32_read_memory_in_3);
  FE_PHC31_read_memory_in_2 : CKBD0BWP7T port map(I => read_memory_in(2), Z => FE_PHN31_read_memory_in_2);
  FE_PHC30_lbl0_booster_sync : DEL0BWP7T port map(I => lbl0_booster_sync, Z => FE_PHN30_lbl0_booster_sync);
  FE_PHC29_read_memory_in_0 : CKBD0BWP7T port map(I => read_memory_in(0), Z => FE_PHN29_read_memory_in_0);
  FE_PHC28_read_memory_in_6 : CKBD0BWP7T port map(I => read_memory_in(6), Z => FE_PHN28_read_memory_in_6);
  FE_PHC27_read_memory_in_1 : CKBD0BWP7T port map(I => read_memory_in(1), Z => FE_PHN27_read_memory_in_1);
  FE_PHC26_lbl2_data_synced_5 : DEL0BWP7T port map(I => lbl2_data_synced(5), Z => FE_PHN26_lbl2_data_synced_5);
  FE_PHC25_lbl2_borders_synced_5 : DEL1BWP7T port map(I => lbl2_borders_synced(5), Z => FE_PHN25_lbl2_borders_synced_5);
  FE_PHC24_lbl2_jumps_synced_3 : DEL1BWP7T port map(I => lbl2_jumps_synced(3), Z => FE_PHN24_lbl2_jumps_synced_3);
  FE_PHC23_lbl2_data_synced_0 : DEL0BWP7T port map(I => lbl2_data_synced(0), Z => FE_PHN23_lbl2_data_synced_0);
  FE_PHC22_lbl2_jumps_synced_7 : DEL1BWP7T port map(I => lbl2_jumps_synced(7), Z => FE_PHN22_lbl2_jumps_synced_7);
  FE_PHC21_lbl2_data_synced_6 : DEL0BWP7T port map(I => lbl2_data_synced(6), Z => FE_PHN21_lbl2_data_synced_6);
  FE_PHC20_lbl2_borders_synced_6 : DEL1BWP7T port map(I => lbl2_borders_synced(6), Z => FE_PHN20_lbl2_borders_synced_6);
  FE_PHC19_lbl2_jumps_synced_5 : DEL1BWP7T port map(I => lbl2_jumps_synced(5), Z => FE_PHN19_lbl2_jumps_synced_5);
  FE_PHC18_lbl2_data_synced_2 : DEL0BWP7T port map(I => lbl2_data_synced(2), Z => FE_PHN18_lbl2_data_synced_2);
  FE_PHC17_lbl2_borders_synced_4 : DEL1BWP7T port map(I => lbl2_borders_synced(4), Z => FE_PHN17_lbl2_borders_synced_4);
  FE_PHC16_lbl2_jumps_synced_4 : DEL1BWP7T port map(I => lbl2_jumps_synced(4), Z => FE_PHN16_lbl2_jumps_synced_4);
  FE_PHC15_lbl2_jumps_synced_2 : DEL1BWP7T port map(I => lbl2_jumps_synced(2), Z => FE_PHN15_lbl2_jumps_synced_2);
  FE_PHC14_lbl2_borders_synced_3 : DEL1BWP7T port map(I => lbl2_borders_synced(3), Z => FE_PHN14_lbl2_borders_synced_3);
  FE_PHC13_lbl2_jumps_synced_0 : DEL1BWP7T port map(I => lbl2_jumps_synced(0), Z => FE_PHN13_lbl2_jumps_synced_0);
  FE_PHC12_lbl2_data_synced_4 : DEL0BWP7T port map(I => lbl2_data_synced(4), Z => FE_PHN12_lbl2_data_synced_4);
  FE_PHC11_lbl2_borders_synced_1 : DEL1BWP7T port map(I => lbl2_borders_synced(1), Z => FE_PHN11_lbl2_borders_synced_1);
  FE_PHC10_lbl2_borders_synced_0 : DEL1BWP7T port map(I => lbl2_borders_synced(0), Z => FE_PHN10_lbl2_borders_synced_0);
  FE_PHC9_lbl2_jumps_synced_6 : DEL1BWP7T port map(I => lbl2_jumps_synced(6), Z => FE_PHN9_lbl2_jumps_synced_6);
  FE_PHC8_lbl2_jumps_synced_1 : DEL1BWP7T port map(I => lbl2_jumps_synced(1), Z => FE_PHN8_lbl2_jumps_synced_1);
  FE_PHC7_lbl2_data_synced_7 : DEL0BWP7T port map(I => lbl2_data_synced(7), Z => FE_PHN7_lbl2_data_synced_7);
  FE_PHC6_lbl2_data_synced_3 : DEL0BWP7T port map(I => lbl2_data_synced(3), Z => FE_PHN6_lbl2_data_synced_3);
  FE_OFC5_memory_enable_out : BUFFD5BWP7T port map(I => FE_OFN5_memory_enable_out, Z => memory_enable_out);
  FE_OFC4_lbl2_n_4 : DEL01BWP7T port map(I => lbl2_n_4, Z => FE_OFN4_lbl2_n_4);
  FE_OFC3_rst : DEL01BWP7T port map(I => rst, Z => FE_OFN3_rst);
  CTS_ccl_a_BUF_clk_G0_L1_2 : CKBD6BWP7T port map(I => clk, Z => CTS_12);
  CTS_ccl_a_BUF_clk_G0_L1_1 : CKBD6BWP7T port map(I => clk, Z => CTS_11);
  FE_DBTC4_rst : INVD2BWP7T port map(I => FE_OFN3_rst, ZN => FE_DBTN4_rst);
  FE_DBTC3_memory_reset_out : CKND1BWP7T port map(I => memory_reset_out, ZN => FE_DBTN3_memory_reset_out);
  FE_DBTC2_lbl2_h_count_3 : INVD1BWP7T port map(I => lbl2_h_count(3), ZN => FE_DBTN2_lbl2_h_count_3);
  FE_DBTC1_lbl2_h_count_1 : INVD0BWP7T port map(I => lbl2_h_count(1), ZN => FE_DBTN1_lbl2_h_count_1);
  FE_DBTC0_lbl2_v_count_2 : INVD1BWP7T port map(I => lbl2_v_count(2), ZN => FE_DBTN0_lbl2_v_count_2);
  lbl2_g2827 : NR4D0BWP7T port map(A1 => lbl2_n_143, A2 => lbl2_n_56, A3 => lbl2_n_125, A4 => lbl2_n_114, ZN => lbl2_n_190);
  lbl2_g2828 : NR4D0BWP7T port map(A1 => lbl2_n_142, A2 => lbl2_n_56, A3 => lbl2_n_126, A4 => lbl2_n_115, ZN => lbl2_n_189);
  lbl2_g2829 : ND4D0BWP7T port map(A1 => lbl2_n_141, A2 => lbl2_n_128, A3 => lbl2_n_121, A4 => lbl2_n_118, ZN => lbl2_n_143);
  lbl2_g2830 : ND4D0BWP7T port map(A1 => lbl2_n_140, A2 => lbl2_n_131, A3 => lbl2_n_119, A4 => lbl2_n_120, ZN => lbl2_n_142);
  lbl2_g2831 : NR3D0BWP7T port map(A1 => lbl2_n_138, A2 => lbl2_n_136, A3 => lbl2_n_129, ZN => lbl2_n_141);
  lbl2_g2832 : NR3D0BWP7T port map(A1 => lbl2_n_139, A2 => lbl2_n_137, A3 => lbl2_n_130, ZN => lbl2_n_140);
  lbl2_g2833 : OAI221D0BWP7T port map(A1 => lbl2_n_123, A2 => position_1(8), B1 => position_1(4), B2 => lbl2_n_124, C => lbl2_n_135, ZN => lbl2_n_139);
  lbl2_g2834 : OAI221D0BWP7T port map(A1 => lbl2_n_123, A2 => position_0(8), B1 => position_0(4), B2 => lbl2_n_124, C => lbl2_n_134, ZN => lbl2_n_138);
  lbl2_g2835 : AO211D0BWP7T port map(A1 => lbl2_n_123, A2 => position_1(8), B => lbl2_n_133, C => lbl2_n_116, Z => lbl2_n_137);
  lbl2_g2836 : AO211D0BWP7T port map(A1 => lbl2_n_123, A2 => position_0(8), B => lbl2_n_132, C => lbl2_n_117, Z => lbl2_n_136);
  lbl2_g2837 : AOI22D0BWP7T port map(A1 => lbl2_n_124, A2 => position_1(4), B1 => lbl2_n_127, B2 => position_1(3), ZN => lbl2_n_135);
  lbl2_g2838 : AOI22D0BWP7T port map(A1 => lbl2_n_124, A2 => position_0(4), B1 => lbl2_n_127, B2 => position_0(3), ZN => lbl2_n_134);
  lbl2_g2839 : NR2D0BWP7T port map(A1 => lbl2_n_127, A2 => position_1(3), ZN => lbl2_n_133);
  lbl2_g2840 : NR2XD0BWP7T port map(A1 => lbl2_n_127, A2 => position_0(3), ZN => lbl2_n_132);
  lbl2_g2841 : XNR2D1BWP7T port map(A1 => lbl2_y_vec(2), A2 => position_1(7), ZN => lbl2_n_131);
  lbl2_g2842 : CKXOR2D1BWP7T port map(A1 => lbl2_y_vec(4), A2 => position_1(9), Z => lbl2_n_130);
  lbl2_g2843 : CKXOR2D1BWP7T port map(A1 => lbl2_y_vec(4), A2 => position_0(9), Z => lbl2_n_129);
  lbl2_g2844 : XNR2D1BWP7T port map(A1 => lbl2_y_vec(2), A2 => position_0(7), ZN => lbl2_n_128);
  lbl2_g2845 : INVD1BWP7T port map(I => lbl2_central_x_vec(7), ZN => lbl2_n_127);
  lbl2_g2846 : MOAI22D1BWP7T port map(A1 => lbl2_n_76, A2 => lbl2_h_count(7), B1 => lbl2_n_76, B2 => lbl2_h_count(7), ZN => lbl2_central_x_vec(7));
  lbl2_g2847 : MAOI22D0BWP7T port map(A1 => lbl2_central_x_vec(6), A2 => position_1(2), B1 => lbl2_central_x_vec(6), B2 => position_1(2), ZN => lbl2_n_126);
  lbl2_g2848 : MAOI22D0BWP7T port map(A1 => lbl2_central_x_vec(6), A2 => position_0(2), B1 => lbl2_central_x_vec(6), B2 => position_0(2), ZN => lbl2_n_125);
  lbl2_g2849 : AO22D0BWP7T port map(A1 => lbl2_n_56, A2 => lbl2_h_count(1), B1 => lbl2_h_count(2), B2 => lbl2_n_156, Z => lbl2_dx(2));
  lbl2_g2850 : AO22D0BWP7T port map(A1 => lbl2_n_56, A2 => lbl2_h_count(2), B1 => lbl2_h_count(3), B2 => lbl2_n_156, Z => lbl2_dx(3));
  lbl2_g2851 : AO22D0BWP7T port map(A1 => lbl2_n_56, A2 => lbl2_v_count(2), B1 => lbl2_v_count(3), B2 => lbl2_n_156, Z => lbl2_dy_vec(3));
  lbl2_g2852 : AO22D0BWP7T port map(A1 => lbl2_n_56, A2 => lbl2_h_count(0), B1 => lbl2_h_count(1), B2 => lbl2_n_156, Z => lbl2_dx(1));
  lbl2_g2853 : AO22D0BWP7T port map(A1 => lbl2_n_56, A2 => lbl2_v_count(1), B1 => lbl2_v_count(2), B2 => lbl2_n_156, Z => lbl2_dy_vec(2));
  lbl2_g2854 : INVD1BWP7T port map(I => lbl2_n_124, ZN => lbl2_central_x_vec(8));
  lbl2_g2856 : AO22D0BWP7T port map(A1 => lbl2_n_56, A2 => lbl2_v_count(0), B1 => lbl2_v_count(1), B2 => lbl2_n_156, Z => lbl2_dy_vec(1));
  lbl2_g2857 : XNR2D1BWP7T port map(A1 => lbl2_n_146, A2 => lbl2_h_count(8), ZN => lbl2_n_124);
  lbl2_g2858 : MOAI22D0BWP7T port map(A1 => lbl2_n_156, A2 => lbl2_v_count(3), B1 => lbl2_n_156, B2 => lbl2_v_count(6), ZN => lbl2_y_vec(2));
  lbl2_g2859 : MOAI22D0BWP7T port map(A1 => lbl2_n_156, A2 => lbl2_v_count(7), B1 => lbl2_n_156, B2 => lbl2_v_count(8), ZN => lbl2_y_vec(4));
  lbl2_g2860 : MAOI22D0BWP7T port map(A1 => lbl2_n_156, A2 => lbl2_v_count(7), B1 => lbl2_n_156, B2 => lbl2_v_count(6), ZN => lbl2_n_123);
  lbl2_g2861 : INR2D1BWP7T port map(A1 => lbl2_v_count(0), B1 => lbl2_n_56, ZN => lbl2_dy_vec(0));
  lbl2_g2862 : CKAN2D1BWP7T port map(A1 => lbl2_n_156, A2 => lbl2_h_count(0), Z => lbl2_dx(0));
  lbl2_g2863 : INVD1BWP7T port map(I => lbl2_n_56, ZN => lbl2_n_156);
  lbl2_g2864 : XNR2D1BWP7T port map(A1 => lbl2_v_count(5), A2 => position_0(6), ZN => lbl2_n_121);
  lbl2_g2865 : XNR2D1BWP7T port map(A1 => lbl2_v_count(4), A2 => position_1(5), ZN => lbl2_n_120);
  lbl2_g2866 : XNR2D1BWP7T port map(A1 => lbl2_v_count(5), A2 => position_1(6), ZN => lbl2_n_119);
  lbl2_g2867 : ND2D1BWP7T port map(A1 => lbl2_n_147, A2 => lbl2_h_count(5), ZN => lbl2_n_146);
  lbl2_g2868 : NR2XD0BWP7T port map(A1 => lbl2_n_158, A2 => game_state(2), ZN => lbl2_n_56);
  lbl2_g2869 : XNR2D1BWP7T port map(A1 => lbl2_v_count(4), A2 => position_0(5), ZN => lbl2_n_118);
  lbl2_g2870 : CKXOR2D1BWP7T port map(A1 => lbl2_h_count(4), A2 => position_0(0), Z => lbl2_n_117);
  lbl2_g2871 : CKXOR2D0BWP7T port map(A1 => lbl2_h_count(4), A2 => position_1(0), Z => lbl2_n_116);
  lbl2_g2872 : MAOI22D0BWP7T port map(A1 => lbl2_central_x_vec(5), A2 => position_1(1), B1 => lbl2_central_x_vec(5), B2 => position_1(1), ZN => lbl2_n_115);
  lbl2_g2873 : MAOI22D0BWP7T port map(A1 => lbl2_central_x_vec(5), A2 => position_0(1), B1 => lbl2_central_x_vec(5), B2 => position_0(1), ZN => lbl2_n_114);
  lbl2_g2874 : MOAI22D1BWP7T port map(A1 => lbl2_central_x_vec(5), A2 => lbl2_h_count(6), B1 => lbl2_central_x_vec(5), B2 => lbl2_h_count(6), ZN => lbl2_central_x_vec(6));
  lbl2_g2875 : AN2D1BWP7T port map(A1 => lbl2_h_count(6), A2 => lbl2_h_count(7), Z => lbl2_n_147);
  lbl2_g2876 : OR2D1BWP7T port map(A1 => game_state(0), A2 => game_state(1), Z => lbl2_n_158);
  lbl2_g2877 : ND2D1BWP7T port map(A1 => lbl2_h_count(5), A2 => lbl2_h_count(6), ZN => lbl2_n_76);
  lbl2_color_reg_0 : DFD0BWP7T port map(CP => CTS_12, D => lbl2_n_104, Q => UNCONNECTED, QN => lbl2_n_109);
  lbl2_color_reg_1 : DFD0BWP7T port map(CP => CTS_12, D => lbl2_n_107, Q => UNCONNECTED0, QN => lbl2_n_111);
  lbl2_color_reg_2 : DFD0BWP7T port map(CP => CTS_12, D => lbl2_n_106, Q => UNCONNECTED1, QN => lbl2_n_112);
  lbl2_color_reg_3 : DFD0BWP7T port map(CP => CTS_12, D => lbl2_n_105, Q => UNCONNECTED2, QN => lbl2_n_110);
  lbl2_h_sync_reg : DFKSND1BWP7T port map(CP => CTS_12, D => lbl2_n_84, Q => UNCONNECTED3, QN => lbl2_n_92, SN => FE_DBTN4_rst);
  lbl2_v_sync_reg : DFKSND0BWP7T port map(CP => CTS_11, D => FE_OFN3_rst, Q => UNCONNECTED4, QN => lbl2_n_101, SN => lbl2_n_94);
  lbl2_g3640 : IINR4D0BWP7T port map(A1 => lbl2_dx(2), A2 => lbl2_dx(3), B1 => lbl2_n_108, B2 => lbl2_n_89, ZN => x_increment);
  lbl2_g3642 : INVD5BWP7T port map(I => lbl2_n_112, ZN => color_out(2));
  lbl2_g3644 : INVD5BWP7T port map(I => lbl2_n_111, ZN => color_out(1));
  lbl2_g3646 : INVD5BWP7T port map(I => lbl2_n_110, ZN => color_out(3));
  lbl2_g3648 : INVD5BWP7T port map(I => lbl2_n_109, ZN => color_out(0));
  lbl2_g3649 : OAI211D1BWP7T port map(A1 => lbl2_n_56, A2 => lbl2_dx(0), B => lbl2_n_103, C => lbl2_dx(1), ZN => lbl2_n_108);
  lbl2_g3650 : AO222D0BWP7T port map(A1 => lbl2_homescreen_color(1), A2 => lbl2_n_99, B1 => lbl2_pixelator_color(1), B2 => lbl2_n_102, C1 => lbl2_sidebar_color(1), C2 => lbl2_n_97, Z => lbl2_n_107);
  lbl2_g3651 : AO222D0BWP7T port map(A1 => lbl2_homescreen_color(2), A2 => lbl2_n_99, B1 => lbl2_pixelator_color(2), B2 => lbl2_n_102, C1 => lbl2_sidebar_color(2), C2 => lbl2_n_97, Z => lbl2_n_106);
  lbl2_g3652 : AO222D0BWP7T port map(A1 => lbl2_homescreen_color(3), A2 => lbl2_n_99, B1 => lbl2_pixelator_color(3), B2 => lbl2_n_102, C1 => lbl2_sidebar_color(3), C2 => lbl2_n_97, Z => lbl2_n_105);
  lbl2_g3653 : AO222D0BWP7T port map(A1 => lbl2_homescreen_color(0), A2 => lbl2_n_99, B1 => lbl2_pixelator_color(0), B2 => lbl2_n_102, C1 => lbl2_sidebar_color(0), C2 => lbl2_n_97, Z => lbl2_n_104);
  lbl2_g3654 : MOAI22D0BWP7T port map(A1 => lbl2_n_100, A2 => lbl2_n_95, B1 => lbl2_n_100, B2 => lbl2_n_95, ZN => lbl2_n_103);
  lbl2_g3655 : INR3D0BWP7T port map(A1 => lbl2_n_70, B1 => lbl2_n_96, B2 => lbl2_n_86, ZN => y_increment);
  lbl2_g3657 : INVD5BWP7T port map(I => lbl2_n_101, ZN => v_sync_out);
  lbl2_g3658 : NR2D1BWP7T port map(A1 => lbl2_n_98, A2 => lbl2_n_56, ZN => lbl2_n_102);
  lbl2_g3659 : INR2XD0BWP7T port map(A1 => lbl2_n_86, B1 => lbl2_n_96, ZN => reset_vga_mem);
  lbl2_g3660 : AOI222D0BWP7T port map(A1 => lbl2_n_56, A2 => lbl2_n_88, B1 => lbl2_n_90, B2 => lbl2_n_74, C1 => lbl2_n_156, C2 => lbl2_h_count(8), ZN => lbl2_n_100);
  lbl2_g3661 : NR2D1BWP7T port map(A1 => lbl2_n_98, A2 => lbl2_n_156, ZN => lbl2_n_99);
  lbl2_g3662 : ND2D1BWP7T port map(A1 => lbl2_n_91, A2 => lbl2_n_93, ZN => lbl2_n_98);
  lbl2_g3663 : INR2D1BWP7T port map(A1 => lbl2_n_93, B1 => lbl2_n_91, ZN => lbl2_n_97);
  lbl2_g3664 : OR4D1BWP7T port map(A1 => lbl2_h_count(3), A2 => lbl2_n_74, A3 => lbl2_n_79, A4 => lbl2_n_89, Z => lbl2_n_96);
  lbl2_g3665 : AO32D1BWP7T port map(A1 => lbl2_n_56, A2 => lbl2_n_87, A3 => lbl2_n_74, B1 => lbl2_n_156, B2 => lbl2_h_count(9), Z => lbl2_n_95);
  lbl2_g3666 : OAI31D0BWP7T port map(A1 => lbl2_v_count(9), A2 => lbl2_v_count(4), A3 => lbl2_n_82, B => FE_DBTN4_rst, ZN => lbl2_n_94);
  lbl2_g3667 : NR4D0BWP7T port map(A1 => lbl2_n_89, A2 => lbl2_n_83, A3 => lbl2_n_80, A4 => FE_OFN3_rst, ZN => lbl2_n_93);
  lbl2_g3669 : INVD5BWP7T port map(I => lbl2_n_92, ZN => h_sync_out);
  lbl2_g3670 : INR3D0BWP7T port map(A1 => lbl2_h_count(6), B1 => lbl2_n_65, B2 => lbl2_n_225, ZN => lbl2_n_90);
  lbl2_g3671 : AOI211XD0BWP7T port map(A1 => lbl2_n_146, A2 => lbl2_n_67, B => lbl2_n_85, C => lbl2_n_69, ZN => lbl2_n_91);
  lbl2_g3672 : OAI21D0BWP7T port map(A1 => lbl2_n_158, A2 => lbl2_n_58, B => busy, ZN => lbl2_n_89);
  lbl2_g3673 : MOAI22D0BWP7T port map(A1 => lbl2_n_76, A2 => lbl2_n_75, B1 => lbl2_n_76, B2 => lbl2_h_count(7), ZN => lbl2_n_88);
  lbl2_g3674 : MOAI22D0BWP7T port map(A1 => lbl2_n_226, A2 => lbl2_h_count(8), B1 => lbl2_n_226, B2 => lbl2_h_count(8), ZN => lbl2_n_87);
  lbl2_g3675 : OAI22D0BWP7T port map(A1 => lbl2_n_71, A2 => lbl2_h_count(5), B1 => lbl2_n_146, B2 => lbl2_n_59, ZN => lbl2_n_85);
  lbl2_g3676 : INR2XD0BWP7T port map(A1 => lbl2_n_78, B1 => lbl2_v_count(9), ZN => busy);
  lbl2_g3677 : NR4D0BWP7T port map(A1 => lbl2_n_227, A2 => lbl2_y_vec(4), A3 => lbl2_v_count(4), A4 => lbl2_v_count(5), ZN => lbl2_n_86);
  lbl2_g3678 : AOI21D0BWP7T port map(A1 => lbl2_n_73, A2 => lbl2_n_76, B => FE_OFN3_rst, ZN => lbl2_n_84);
  lbl2_g3679 : OA21D0BWP7T port map(A1 => lbl2_n_72, A2 => lbl2_n_75, B => lbl2_n_69, Z => lbl2_n_83);
  lbl2_g3680 : IIND4D0BWP7T port map(A1 => lbl2_n_78, A2 => lbl2_v_count(2), B1 => lbl2_v_count(3), B2 => lbl2_v_count(1), ZN => lbl2_n_82);
  lbl2_g3682 : AOI211XD0BWP7T port map(A1 => lbl2_n_148, A2 => lbl2_h_count(7), B => lbl2_n_147, C => lbl2_n_68, ZN => lbl2_n_80);
  lbl2_g3683 : OR4D1BWP7T port map(A1 => lbl2_h_count(1), A2 => lbl2_h_count(2), A3 => lbl2_h_count(0), A4 => lbl2_n_72, Z => lbl2_n_79);
  lbl2_g3684 : ND4D0BWP7T port map(A1 => lbl2_v_count(5), A2 => lbl2_v_count(7), A3 => lbl2_v_count(8), A4 => lbl2_v_count(6), ZN => lbl2_n_78);
  lbl2_g3687 : INVD1BWP7T port map(I => lbl2_n_73, ZN => lbl2_n_74);
  lbl2_g3688 : IND2D1BWP7T port map(A1 => lbl2_h_count(7), B1 => lbl2_n_68, ZN => lbl2_n_75);
  lbl2_g3689 : NR2XD0BWP7T port map(A1 => lbl2_n_68, A2 => lbl2_h_count(7), ZN => lbl2_n_73);
  lbl2_g3690 : ND3D0BWP7T port map(A1 => lbl2_central_x_vec(8), A2 => lbl2_central_x_vec(7), A3 => lbl2_central_x_vec(6), ZN => lbl2_n_71);
  lbl2_g3691 : NR4D0BWP7T port map(A1 => lbl2_dy_vec(1), A2 => lbl2_dy_vec(2), A3 => lbl2_dy_vec(3), A4 => lbl2_dy_vec(0), ZN => lbl2_n_70);
  lbl2_g3692 : IND2D1BWP7T port map(A1 => lbl2_h_count(6), B1 => lbl2_n_65, ZN => lbl2_n_72);
  lbl2_g3693 : INVD1BWP7T port map(I => lbl2_n_67, ZN => lbl2_n_68);
  lbl2_g3694 : ND2D0BWP7T port map(A1 => lbl2_h_count(5), A2 => lbl2_h_count(3), ZN => lbl2_n_66);
  lbl2_g3695 : CKAN2D1BWP7T port map(A1 => lbl2_h_count(9), A2 => lbl2_h_count(8), Z => lbl2_n_69);
  lbl2_g3696 : NR2XD0BWP7T port map(A1 => lbl2_h_count(9), A2 => lbl2_h_count(8), ZN => lbl2_n_67);
  lbl2_g3699 : NR2XD0BWP7T port map(A1 => lbl2_h_count(5), A2 => lbl2_h_count(4), ZN => lbl2_n_65);
  lbl2_g3704 : CKND1BWP7T port map(I => game_state(2), ZN => lbl2_n_58);
  lbl2_g2126 : MOAI22D0BWP7T port map(A1 => lbl2_n_52, A2 => lbl2_h_count(5), B1 => lbl2_n_52, B2 => lbl2_h_count(5), ZN => lbl2_n_150);
  lbl2_g2127 : MOAI22D1BWP7T port map(A1 => lbl2_n_53, A2 => lbl2_h_count(6), B1 => lbl2_n_53, B2 => lbl2_h_count(6), ZN => lbl2_n_151);
  lbl2_g2128 : IOA21D1BWP7T port map(A1 => lbl2_h_count(4), A2 => lbl2_h_count(9), B => lbl2_n_52, ZN => lbl2_n_149);
  lbl2_g2129 : INR2D1BWP7T port map(A1 => lbl2_n_148, B1 => lbl2_h_count(9), ZN => lbl2_n_53);
  lbl2_g2130 : CKMUX2D1BWP7T port map(I0 => player_state_0(0), I1 => player_state_1(0), S => lbl2_h_count(9), Z => lbl2_n_152);
  lbl2_g2131 : MUX2D1BWP7T port map(I0 => direction_in(1), I1 => direction_in(3), S => lbl2_h_count(9), Z => lbl2_n_154);
  lbl2_g2132 : MUX2D1BWP7T port map(I0 => direction_in(0), I1 => direction_in(2), S => lbl2_h_count(9), Z => lbl2_n_153);
  lbl2_g2133 : OR2D1BWP7T port map(A1 => lbl2_h_count(5), A2 => lbl2_h_count(4), Z => lbl2_n_148);
  lbl2_g2134 : OR2D1BWP7T port map(A1 => lbl2_h_count(4), A2 => lbl2_h_count(9), Z => lbl2_n_52);
  lbl2_borders_synced_reg_0 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN10_lbl2_borders_synced_0, DB => borders(0), Q => lbl2_borders_synced(0), SA => FE_OFN4_lbl2_n_4);
  lbl2_borders_synced_reg_1 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN11_lbl2_borders_synced_1, DB => borders(1), Q => lbl2_borders_synced(1), SA => FE_OFN4_lbl2_n_4);
  lbl2_borders_synced_reg_2 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN41_lbl2_borders_synced_2, DB => borders(2), Q => lbl2_borders_synced(2), SA => FE_OFN4_lbl2_n_4);
  lbl2_borders_synced_reg_3 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN14_lbl2_borders_synced_3, DB => borders(3), Q => lbl2_borders_synced(3), SA => FE_OFN4_lbl2_n_4);
  lbl2_borders_synced_reg_4 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN17_lbl2_borders_synced_4, DB => borders(4), Q => lbl2_borders_synced(4), SA => FE_OFN4_lbl2_n_4);
  lbl2_borders_synced_reg_5 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN25_lbl2_borders_synced_5, DB => borders(5), Q => lbl2_borders_synced(5), SA => FE_OFN4_lbl2_n_4);
  lbl2_borders_synced_reg_6 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN20_lbl2_borders_synced_6, DB => borders(6), Q => lbl2_borders_synced(6), SA => FE_OFN4_lbl2_n_4);
  lbl2_borders_synced_reg_7 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN35_lbl2_borders_synced_7, DB => borders(7), Q => lbl2_borders_synced(7), SA => FE_OFN4_lbl2_n_4);
  lbl2_data_synced_reg_0 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN23_lbl2_data_synced_0, DB => FE_PHN29_read_memory_in_0, Q => lbl2_data_synced(0), SA => FE_OFN4_lbl2_n_4);
  lbl2_data_synced_reg_1 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN38_lbl2_data_synced_1, DB => FE_PHN27_read_memory_in_1, Q => lbl2_data_synced(1), SA => FE_OFN4_lbl2_n_4);
  lbl2_data_synced_reg_2 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN18_lbl2_data_synced_2, DB => FE_PHN31_read_memory_in_2, Q => lbl2_data_synced(2), SA => FE_OFN4_lbl2_n_4);
  lbl2_data_synced_reg_3 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN6_lbl2_data_synced_3, DB => FE_PHN32_read_memory_in_3, Q => lbl2_data_synced(3), SA => FE_OFN4_lbl2_n_4);
  lbl2_data_synced_reg_4 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN12_lbl2_data_synced_4, DB => FE_PHN34_read_memory_in_4, Q => lbl2_data_synced(4), SA => FE_OFN4_lbl2_n_4);
  lbl2_data_synced_reg_5 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN26_lbl2_data_synced_5, DB => FE_PHN33_read_memory_in_5, Q => lbl2_data_synced(5), SA => FE_OFN4_lbl2_n_4);
  lbl2_data_synced_reg_6 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN21_lbl2_data_synced_6, DB => FE_PHN28_read_memory_in_6, Q => lbl2_data_synced(6), SA => FE_OFN4_lbl2_n_4);
  lbl2_data_synced_reg_7 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN7_lbl2_data_synced_7, DB => FE_PHN64_read_memory_in_7, Q => lbl2_data_synced(7), SA => FE_OFN4_lbl2_n_4);
  lbl2_h_count_reg_0 : DFKCNQD1BWP7T port map(CN => lbl2_n_23, CP => CTS_11, D => lbl2_n_11, Q => lbl2_h_count(0));
  lbl2_h_count_reg_1 : DFKCNQD1BWP7T port map(CN => lbl2_n_11, CP => CTS_11, D => lbl2_n_27, Q => lbl2_h_count(1));
  lbl2_h_count_reg_2 : DFKCNQD1BWP7T port map(CN => lbl2_n_11, CP => CTS_11, D => lbl2_n_30, Q => lbl2_h_count(2));
  lbl2_h_count_reg_3 : DFKCNQD1BWP7T port map(CN => lbl2_n_11, CP => CTS_11, D => lbl2_n_33, Q => lbl2_h_count(3));
  lbl2_h_count_reg_4 : DFKCNQD1BWP7T port map(CN => lbl2_n_11, CP => CTS_11, D => lbl2_n_36, Q => lbl2_h_count(4));
  lbl2_h_count_reg_6 : DFKCNQD1BWP7T port map(CN => lbl2_n_11, CP => CTS_11, D => lbl2_n_42, Q => lbl2_h_count(6));
  lbl2_h_count_reg_7 : DFKCNQD1BWP7T port map(CN => lbl2_n_11, CP => CTS_11, D => lbl2_n_45, Q => lbl2_h_count(7));
  lbl2_h_count_reg_8 : DFKCNQD1BWP7T port map(CN => lbl2_n_11, CP => CTS_11, D => lbl2_n_48, Q => lbl2_h_count(8));
  lbl2_jumps_synced_reg_0 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN13_lbl2_jumps_synced_0, DB => ramps(0), Q => lbl2_jumps_synced(0), SA => FE_OFN4_lbl2_n_4);
  lbl2_jumps_synced_reg_1 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN8_lbl2_jumps_synced_1, DB => ramps(1), Q => lbl2_jumps_synced(1), SA => FE_OFN4_lbl2_n_4);
  lbl2_jumps_synced_reg_2 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN15_lbl2_jumps_synced_2, DB => ramps(2), Q => lbl2_jumps_synced(2), SA => FE_OFN4_lbl2_n_4);
  lbl2_jumps_synced_reg_3 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN24_lbl2_jumps_synced_3, DB => ramps(3), Q => lbl2_jumps_synced(3), SA => FE_OFN4_lbl2_n_4);
  lbl2_jumps_synced_reg_4 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN16_lbl2_jumps_synced_4, DB => ramps(4), Q => lbl2_jumps_synced(4), SA => FE_OFN4_lbl2_n_4);
  lbl2_jumps_synced_reg_5 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN19_lbl2_jumps_synced_5, DB => ramps(5), Q => lbl2_jumps_synced(5), SA => FE_OFN4_lbl2_n_4);
  lbl2_jumps_synced_reg_6 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN9_lbl2_jumps_synced_6, DB => ramps(6), Q => lbl2_jumps_synced(6), SA => FE_OFN4_lbl2_n_4);
  lbl2_jumps_synced_reg_7 : DFXQD1BWP7T port map(CP => CTS_12, DA => FE_PHN22_lbl2_jumps_synced_7, DB => ramps(7), Q => lbl2_jumps_synced(7), SA => FE_OFN4_lbl2_n_4);
  lbl2_v_count_reg_0 : DFQD1BWP7T port map(CP => CTS_11, D => lbl2_n_25, Q => lbl2_v_count(0));
  lbl2_v_count_reg_1 : DFQD1BWP7T port map(CP => CTS_11, D => lbl2_n_28, Q => lbl2_v_count(1));
  lbl2_v_count_reg_2 : DFQD1BWP7T port map(CP => CTS_11, D => lbl2_n_31, Q => lbl2_v_count(2));
  lbl2_v_count_reg_3 : DFQD1BWP7T port map(CP => CTS_11, D => lbl2_n_34, Q => lbl2_v_count(3));
  lbl2_v_count_reg_4 : DFQD1BWP7T port map(CP => CTS_11, D => lbl2_n_37, Q => lbl2_v_count(4));
  lbl2_v_count_reg_5 : DFQD1BWP7T port map(CP => CTS_11, D => lbl2_n_40, Q => lbl2_v_count(5));
  lbl2_v_count_reg_6 : DFQD1BWP7T port map(CP => CTS_11, D => lbl2_n_43, Q => lbl2_v_count(6));
  lbl2_v_count_reg_7 : DFQD1BWP7T port map(CP => CTS_11, D => lbl2_n_46, Q => lbl2_v_count(7));
  lbl2_v_count_reg_8 : DFQD1BWP7T port map(CP => CTS_11, D => lbl2_n_49, Q => lbl2_v_count(8));
  lbl2_v_count_reg_9 : DFQD1BWP7T port map(CP => CTS_11, D => lbl2_n_51, Q => FE_PHN63_lbl2_v_count_9);
  lbl2_g3244 : AO22D0BWP7T port map(A1 => lbl2_n_50, A2 => lbl2_n_22, B1 => lbl2_v_count(9), B2 => lbl2_n_11, Z => lbl2_n_51);
  lbl2_g3247 : AO22D0BWP7T port map(A1 => lbl2_n_48, A2 => lbl2_n_22, B1 => FE_PHN44_lbl2_v_count_8, B2 => lbl2_n_11, Z => lbl2_n_49);
  lbl2_g3248 : MOAI22D0BWP7T port map(A1 => lbl2_n_47, A2 => lbl2_n_17, B1 => lbl2_n_47, B2 => lbl2_n_17, ZN => lbl2_n_50);
  lbl2_g3249 : HA1D0BWP7T port map(A => lbl2_n_13, B => lbl2_n_44, CO => lbl2_n_47, S => lbl2_n_48);
  lbl2_g3252 : AO22D0BWP7T port map(A1 => lbl2_n_45, A2 => lbl2_n_22, B1 => FE_PHN45_lbl2_v_count_7, B2 => lbl2_n_11, Z => lbl2_n_46);
  lbl2_g3253 : HA1D0BWP7T port map(A => lbl2_n_18, B => lbl2_n_41, CO => lbl2_n_44, S => lbl2_n_45);
  lbl2_g3256 : AO22D0BWP7T port map(A1 => lbl2_n_42, A2 => lbl2_n_22, B1 => FE_PHN52_lbl2_v_count_6, B2 => lbl2_n_11, Z => lbl2_n_43);
  lbl2_g3257 : HA1D0BWP7T port map(A => lbl2_n_20, B => lbl2_n_38, CO => lbl2_n_41, S => lbl2_n_42);
  lbl2_g3260 : AO22D0BWP7T port map(A1 => lbl2_n_39, A2 => lbl2_n_22, B1 => lbl2_v_count(5), B2 => lbl2_n_11, Z => lbl2_n_40);
  lbl2_g3261 : HA1D0BWP7T port map(A => lbl2_n_19, B => lbl2_n_35, CO => lbl2_n_38, S => lbl2_n_39);
  lbl2_g3264 : AO22D0BWP7T port map(A1 => lbl2_n_36, A2 => lbl2_n_22, B1 => lbl2_v_count(4), B2 => lbl2_n_11, Z => lbl2_n_37);
  lbl2_g3265 : HA1D0BWP7T port map(A => lbl2_n_14, B => lbl2_n_32, CO => lbl2_n_35, S => lbl2_n_36);
  lbl2_g3268 : AO22D0BWP7T port map(A1 => lbl2_n_33, A2 => lbl2_n_22, B1 => lbl2_v_count(3), B2 => lbl2_n_11, Z => lbl2_n_34);
  lbl2_g3269 : HA1D0BWP7T port map(A => lbl2_n_15, B => lbl2_n_29, CO => lbl2_n_32, S => lbl2_n_33);
  lbl2_g3272 : AO22D0BWP7T port map(A1 => lbl2_n_30, A2 => lbl2_n_22, B1 => lbl2_v_count(2), B2 => lbl2_n_11, Z => lbl2_n_31);
  lbl2_g3273 : HA1D0BWP7T port map(A => lbl2_n_16, B => lbl2_n_26, CO => lbl2_n_29, S => lbl2_n_30);
  lbl2_g3276 : AO22D0BWP7T port map(A1 => lbl2_n_27, A2 => lbl2_n_22, B1 => lbl2_v_count(1), B2 => lbl2_n_11, Z => lbl2_n_28);
  lbl2_g3277 : HA1D0BWP7T port map(A => lbl2_n_24, B => lbl2_n_12, CO => lbl2_n_26, S => lbl2_n_27);
  lbl2_g3280 : MOAI22D0BWP7T port map(A1 => lbl2_n_21, A2 => lbl2_n_24, B1 => lbl2_n_11, B2 => lbl2_v_count(0), ZN => lbl2_n_25);
  lbl2_g3281 : INVD0BWP7T port map(I => lbl2_n_23, ZN => lbl2_n_24);
  lbl2_g3282 : INVD0BWP7T port map(I => lbl2_n_22, ZN => lbl2_n_21);
  lbl2_g3283 : AO21D0BWP7T port map(A1 => lbl2_n_9, A2 => lbl2_v_count(6), B => lbl2_h_count(6), Z => lbl2_n_20);
  lbl2_g3284 : AO21D0BWP7T port map(A1 => lbl2_n_9, A2 => lbl2_v_count(5), B => lbl2_h_count(5), Z => lbl2_n_19);
  lbl2_g3285 : AO21D0BWP7T port map(A1 => lbl2_n_9, A2 => lbl2_v_count(7), B => lbl2_h_count(7), Z => lbl2_n_18);
  lbl2_g3286 : AOI22D0BWP7T port map(A1 => lbl2_n_9, A2 => lbl2_v_count(0), B1 => lbl2_n_10, B2 => lbl2_h_count(0), ZN => lbl2_n_23);
  lbl2_g3287 : AOI211XD0BWP7T port map(A1 => lbl2_n_8, A2 => lbl2_v_count(9), B => lbl2_n_10, C => FE_OFN3_rst, ZN => lbl2_n_22);
  lbl2_g3288 : AOI22D0BWP7T port map(A1 => lbl2_n_9, A2 => lbl2_v_count(9), B1 => lbl2_n_10, B2 => lbl2_h_count(9), ZN => lbl2_n_17);
  lbl2_g3289 : AO22D0BWP7T port map(A1 => lbl2_n_9, A2 => lbl2_v_count(2), B1 => lbl2_h_count(2), B2 => lbl2_n_10, Z => lbl2_n_16);
  lbl2_g3290 : AO22D0BWP7T port map(A1 => lbl2_n_9, A2 => lbl2_v_count(3), B1 => lbl2_h_count(3), B2 => lbl2_n_10, Z => lbl2_n_15);
  lbl2_g3291 : AO22D0BWP7T port map(A1 => lbl2_n_9, A2 => lbl2_v_count(4), B1 => lbl2_h_count(4), B2 => lbl2_n_10, Z => lbl2_n_14);
  lbl2_g3292 : AO22D0BWP7T port map(A1 => lbl2_n_9, A2 => lbl2_v_count(8), B1 => lbl2_h_count(8), B2 => lbl2_n_10, Z => lbl2_n_13);
  lbl2_g3293 : AO22D0BWP7T port map(A1 => lbl2_n_9, A2 => lbl2_v_count(1), B1 => lbl2_h_count(1), B2 => lbl2_n_10, Z => lbl2_n_12);
  lbl2_g3294 : NR2XD0BWP7T port map(A1 => lbl2_n_9, A2 => FE_OFN3_rst, ZN => lbl2_n_11);
  lbl2_g3295 : INVD1BWP7T port map(I => lbl2_n_10, ZN => lbl2_n_9);
  lbl2_g3296 : IND4D0BWP7T port map(A1 => lbl2_h_count(7), B1 => lbl2_h_count(8), B2 => lbl2_h_count(9), B3 => lbl2_n_7, ZN => lbl2_n_10);
  lbl2_g3297 : INR4D0BWP7T port map(A1 => lbl2_n_6, B1 => lbl2_v_count(8), B2 => lbl2_v_count(7), B3 => lbl2_v_count(6), ZN => lbl2_n_8);
  lbl2_g3310 : INR4D0BWP7T port map(A1 => lbl2_h_count(4), B1 => lbl2_h_count(6), B2 => lbl2_h_count(5), B3 => lbl2_n_3, ZN => lbl2_n_7);
  lbl2_g3323 : NR3D0BWP7T port map(A1 => lbl2_n_5, A2 => lbl2_v_count(5), A3 => lbl2_v_count(4), ZN => lbl2_n_6);
  lbl2_g3324 : IIND4D0BWP7T port map(A1 => lbl2_v_count(0), A2 => lbl2_v_count(1), B1 => lbl2_v_count(2), B2 => lbl2_v_count(3), ZN => lbl2_n_5);
  lbl2_g3325 : ND4D0BWP7T port map(A1 => lbl2_h_count(0), A2 => lbl2_h_count(2), A3 => lbl2_h_count(1), A4 => lbl2_h_count(3), ZN => lbl2_n_3);
  lbl2_g3326 : ND4D0BWP7T port map(A1 => lbl2_n_2, A2 => lbl2_dx(1), A3 => lbl2_dx(3), A4 => lbl2_dx(2), ZN => lbl2_n_4);
  lbl2_g3327 : IND2D1BWP7T port map(A1 => lbl2_dx(0), B1 => lbl2_n_156, ZN => lbl2_n_2);
  lbl2_g2 : AOI22D0BWP7T port map(A1 => lbl2_n_56, A2 => lbl2_n_66, B1 => lbl2_n_156, B2 => lbl2_h_count(7), ZN => lbl2_n_225);
  lbl2_g3713 : INR2D1BWP7T port map(A1 => lbl2_h_count(3), B1 => lbl2_n_146, ZN => lbl2_n_226);
  lbl2_h_count_reg_5 : DFKCND1BWP7T port map(CN => lbl2_n_11, CP => CTS_11, D => lbl2_n_39, Q => lbl2_h_count(5), QN => lbl2_central_x_vec(5));
  lbl2_h_count_reg_9 : DFKCND1BWP7T port map(CN => lbl2_n_11, CP => CTS_11, D => lbl2_n_50, Q => lbl2_h_count(9), QN => lbl2_n_59);
  lbl2_g3718 : IND2D1BWP7T port map(A1 => lbl2_y_vec(2), B1 => lbl2_n_123, ZN => lbl2_n_227);
  lbl2_dec0_g100 : AO22D0BWP7T port map(A1 => lbl2_dec0_n_2, A2 => lbl2_data_synced(0), B1 => lbl2_data_synced(1), B2 => lbl2_dec0_n_1, Z => lbl2_walls(2));
  lbl2_dec0_g101 : IOA21D1BWP7T port map(A1 => lbl2_dec0_n_2, A2 => lbl2_dec0_n_0, B => lbl2_dec0_n_5, ZN => lbl2_walls(0));
  lbl2_dec0_g102 : IND2D1BWP7T port map(A1 => lbl2_dec0_n_2, B1 => lbl2_dec0_n_3, ZN => lbl2_walls(1));
  lbl2_dec0_g103 : IOA21D1BWP7T port map(A1 => lbl2_dec0_n_0, A2 => lbl2_data_synced(2), B => lbl2_data_synced(1), ZN => lbl2_dec0_n_5);
  lbl2_dec0_g104 : IOA21D1BWP7T port map(A1 => lbl2_data_synced(1), A2 => lbl2_data_synced(2), B => lbl2_dec0_n_3, ZN => lbl2_walls(3));
  lbl2_dec0_g105 : IND2D1BWP7T port map(A1 => lbl2_data_synced(2), B1 => lbl2_data_synced(0), ZN => lbl2_dec0_n_3);
  lbl2_dec0_g106 : ND2D0BWP7T port map(A1 => lbl2_data_synced(0), A2 => lbl2_data_synced(2), ZN => lbl2_dec0_n_1);
  lbl2_dec0_g107 : INR2D1BWP7T port map(A1 => lbl2_data_synced(2), B1 => lbl2_data_synced(1), ZN => lbl2_dec0_n_2);
  lbl2_dec0_g108 : CKND1BWP7T port map(I => lbl2_data_synced(0), ZN => lbl2_dec0_n_0);
  lbl4_g7865 : ND2D1BWP7T port map(A1 => lbl4_n_142, A2 => lbl4_n_66, ZN => borders(6));
  lbl4_g7866 : IND3D1BWP7T port map(A1 => ramps(0), B1 => lbl4_n_84, B2 => lbl4_n_138, ZN => borders(4));
  lbl4_g7867 : IND3D1BWP7T port map(A1 => ramps(7), B1 => lbl4_n_113, B2 => lbl4_n_134, ZN => borders(3));
  lbl4_g7868 : IND2D1BWP7T port map(A1 => ramps(5), B1 => lbl4_n_139, ZN => borders(1));
  lbl4_g7869 : IND3D1BWP7T port map(A1 => ramps(4), B1 => lbl4_n_84, B2 => lbl4_n_131, ZN => borders(0));
  lbl4_g7870 : IND4D0BWP7T port map(A1 => ramps(6), B1 => lbl4_n_66, B2 => lbl4_n_97, B3 => lbl4_n_122, ZN => borders(2));
  lbl4_g7871 : AOI211XD0BWP7T port map(A1 => lbl4_n_127, A2 => lbl4_n_29, B => ramps(2), C => lbl4_n_91, ZN => lbl4_n_142);
  lbl4_g7872 : IND4D0BWP7T port map(A1 => lbl4_n_125, B1 => lbl4_n_106, B2 => lbl4_n_121, B3 => lbl4_n_124, ZN => borders(7));
  lbl4_g7873 : ND3D0BWP7T port map(A1 => lbl4_n_132, A2 => lbl4_n_123, A3 => lbl4_n_116, ZN => borders(5));
  lbl4_g7874 : AOI211XD0BWP7T port map(A1 => lbl4_n_42, A2 => lbl4_n_35, B => lbl4_n_129, C => lbl4_n_102, ZN => lbl4_n_139);
  lbl4_g7875 : AOI22D0BWP7T port map(A1 => lbl4_n_127, A2 => lbl4_n_11, B1 => lbl4_n_92, B2 => lbl4_n_44, ZN => lbl4_n_138);
  lbl4_g7876 : OAI21D0BWP7T port map(A1 => lbl4_n_95, A2 => lbl4_n_20, B => lbl4_n_124, ZN => ramps(3));
  lbl4_g7877 : AOI31D0BWP7T port map(A1 => lbl4_n_3, A2 => lbl4_n_107, A3 => lbl4_n_4, B => lbl4_n_110, ZN => lbl4_n_134);
  lbl4_g7878 : OAI221D0BWP7T port map(A1 => lbl4_n_95, A2 => lbl4_n_14, B1 => lbl4_n_33, B2 => lbl4_n_104, C => lbl4_n_115, ZN => ramps(5));
  lbl4_g7879 : OAI31D1BWP7T port map(A1 => lbl4_n_33, A2 => lbl4_n_58, A3 => lbl4_n_80, B => lbl4_n_126, ZN => ramps(7));
  lbl4_g7880 : AOI33D1BWP7T port map(A1 => lbl4_n_3, A2 => lbl4_n_161, A3 => x_address(0), B1 => start_position_0(3), B2 => lbl4_n_100, B3 => lbl4_n_78, ZN => lbl4_n_132);
  lbl4_g7881 : AOI22D0BWP7T port map(A1 => lbl4_n_118, A2 => lbl4_n_11, B1 => lbl4_n_92, B2 => lbl4_n_74, ZN => lbl4_n_131);
  lbl4_g7882 : OAI31D0BWP7T port map(A1 => lbl4_n_17, A2 => lbl4_n_43, A3 => lbl4_n_80, B => lbl4_n_123, ZN => ramps(1));
  lbl4_g7883 : AO33D0BWP7T port map(A1 => lbl4_n_3, A2 => lbl4_n_107, A3 => x_address(0), B1 => start_position_0(3), B2 => lbl4_n_99, B3 => lbl4_n_78, Z => lbl4_n_129);
  lbl4_g7884 : OAI33D1BWP7T port map(A1 => lbl4_n_21, A2 => lbl4_n_15, A3 => lbl4_n_111, B1 => lbl4_n_49, B2 => lbl4_n_41, B3 => lbl4_n_65, ZN => ramps(2));
  lbl4_g7885 : AOI32D1BWP7T port map(A1 => lbl4_n_103, A2 => lbl4_n_70, A3 => x_address(0), B1 => lbl4_n_89, B2 => lbl4_n_13, ZN => lbl4_n_126);
  lbl4_g7886 : AN3D0BWP7T port map(A1 => lbl4_n_3, A2 => lbl4_n_161, A3 => lbl4_n_4, Z => lbl4_n_125);
  lbl4_g7887 : OAI32D1BWP7T port map(A1 => lbl4_n_12, A2 => lbl4_n_64, A3 => lbl4_n_65, B1 => lbl4_n_61, B2 => lbl4_n_111, ZN => ramps(4));
  lbl4_g7888 : OAI31D0BWP7T port map(A1 => y_address(2), A2 => lbl4_n_47, A3 => lbl4_n_81, B => lbl4_n_117, ZN => lbl4_n_127);
  lbl4_g7889 : AOI22D0BWP7T port map(A1 => lbl4_n_112, A2 => lbl4_n_29, B1 => lbl4_n_105, B2 => lbl4_n_40, ZN => lbl4_n_122);
  lbl4_g7890 : MAOI22D0BWP7T port map(A1 => lbl4_n_100, A2 => lbl4_n_98, B1 => lbl4_n_109, B2 => lbl4_n_20, ZN => lbl4_n_121);
  lbl4_g7891 : IAO21D0BWP7T port map(A1 => lbl4_n_104, A2 => lbl4_n_14, B => lbl4_n_114, ZN => lbl4_n_124);
  lbl4_g7892 : AOI32D1BWP7T port map(A1 => lbl4_n_103, A2 => lbl4_n_57, A3 => lbl4_n_13, B1 => lbl4_n_89, B2 => lbl4_n_34, ZN => lbl4_n_123);
  lbl4_g7893 : AO21D0BWP7T port map(A1 => lbl4_n_105, A2 => lbl4_n_5, B => lbl4_n_112, Z => lbl4_n_118);
  lbl4_g7894 : OA31D1BWP7T port map(A1 => lbl4_n_32, A2 => lbl4_n_15, A3 => lbl4_n_87, B => lbl4_n_90, Z => lbl4_n_117);
  lbl4_g7895 : INR2D1BWP7T port map(A1 => lbl4_n_108, B1 => lbl4_n_21, ZN => ramps(6));
  lbl4_g7896 : INR2D1BWP7T port map(A1 => lbl4_n_108, B1 => lbl4_n_23, ZN => ramps(0));
  lbl4_g7897 : OA32D1BWP7T port map(A1 => lbl4_n_29, A2 => lbl4_n_64, A3 => lbl4_n_75, B1 => lbl4_n_43, B2 => lbl4_n_101, Z => lbl4_n_116);
  lbl4_g7898 : IND3D1BWP7T port map(A1 => lbl4_n_36, B1 => lbl4_n_42, B2 => lbl4_n_103, ZN => lbl4_n_115);
  lbl4_g7899 : AN3D0BWP7T port map(A1 => lbl4_n_103, A2 => lbl4_n_51, A3 => lbl4_n_34, Z => lbl4_n_114);
  lbl4_g7900 : MAOI22D0BWP7T port map(A1 => lbl4_n_99, A2 => lbl4_n_98, B1 => lbl4_n_55, B2 => lbl4_n_20, ZN => lbl4_n_113);
  lbl4_g7901 : NR4D0BWP7T port map(A1 => lbl4_n_77, A2 => lbl4_n_83, A3 => lbl4_n_22, A4 => lbl4_n_4, ZN => lbl4_n_110);
  lbl4_g7902 : CKAN2D1BWP7T port map(A1 => lbl4_n_96, A2 => lbl4_n_55, Z => lbl4_n_109);
  lbl4_g7903 : MOAI22D0BWP7T port map(A1 => lbl4_n_86, A2 => lbl4_n_15, B1 => lbl4_n_82, B2 => lbl4_n_44, ZN => lbl4_n_112);
  lbl4_g7904 : AOI31D0BWP7T port map(A1 => lbl4_n_3, A2 => lbl4_n_73, A3 => lbl4_n_25, B => lbl4_n_93, ZN => lbl4_n_111);
  lbl4_g7905 : OR4XD1BWP7T port map(A1 => lbl4_n_4, A2 => lbl4_n_29, A3 => lbl4_n_64, A4 => lbl4_n_83, Z => lbl4_n_106);
  lbl4_g7906 : OAI32D1BWP7T port map(A1 => lbl4_n_26, A2 => lbl4_n_79, A3 => map_selected(1), B1 => lbl4_n_38, B2 => lbl4_n_94, ZN => lbl4_n_108);
  lbl4_g7908 : AO32D1BWP7T port map(A1 => lbl4_n_63, A2 => lbl4_n_54, A3 => lbl4_n_25, B1 => lbl4_n_88, B2 => lbl4_n_70, Z => lbl4_n_107);
  lbl4_g7909 : NR3D0BWP7T port map(A1 => lbl4_n_77, A2 => lbl4_n_75, A3 => lbl4_n_22, ZN => lbl4_n_102);
  lbl4_g7910 : IAO21D0BWP7T port map(A1 => lbl4_n_80, A2 => x_address(4), B => lbl4_n_35, ZN => lbl4_n_101);
  lbl4_g7911 : NR2D1BWP7T port map(A1 => lbl4_n_87, A2 => lbl4_n_52, ZN => lbl4_n_105);
  lbl4_g7912 : IND4D0BWP7T port map(A1 => lbl4_n_32, B1 => lbl4_n_6, B2 => lbl4_n_59, B3 => lbl4_n_69, ZN => lbl4_n_104);
  lbl4_g7913 : AOI211D1BWP7T port map(A1 => lbl4_n_71, A2 => y_address(4), B => lbl4_n_27, C => lbl4_n_72, ZN => lbl4_n_103);
  lbl4_g7914 : ND3D0BWP7T port map(A1 => lbl4_n_74, A2 => lbl4_n_68, A3 => lbl4_n_11, ZN => lbl4_n_97);
  lbl4_g7915 : IND3D0BWP7T port map(A1 => lbl4_n_80, B1 => x_address(4), B2 => x_address(2), ZN => lbl4_n_96);
  lbl4_g7916 : OAI32D0BWP7T port map(A1 => y_address(3), A2 => lbl4_n_38, A3 => lbl4_n_46, B1 => y_address(4), B2 => lbl4_n_76, ZN => lbl4_n_100);
  lbl4_g7917 : MOAI22D0BWP7T port map(A1 => lbl4_n_76, A2 => lbl4_n_6, B1 => lbl4_n_63, B2 => lbl4_n_8, ZN => lbl4_n_99);
  lbl4_g7918 : AOI211D1BWP7T port map(A1 => lbl4_n_67, A2 => lbl4_n_45, B => lbl4_n_27, C => lbl4_n_4, ZN => lbl4_n_98);
  lbl4_g7919 : CKND1BWP7T port map(I => lbl4_n_93, ZN => lbl4_n_94);
  lbl4_g7920 : AN3D0BWP7T port map(A1 => lbl4_n_68, A2 => lbl4_n_44, A3 => lbl4_n_11, Z => lbl4_n_91);
  lbl4_g7921 : OAI21D0BWP7T port map(A1 => lbl4_n_70, A2 => lbl4_n_54, B => lbl4_n_82, ZN => lbl4_n_90);
  lbl4_g7922 : IND2D1BWP7T port map(A1 => lbl4_n_80, B1 => lbl4_n_51, ZN => lbl4_n_95);
  lbl4_g7923 : AOI211D1BWP7T port map(A1 => lbl4_n_56, A2 => lbl4_n_45, B => lbl4_n_27, C => y_address(3), ZN => lbl4_n_93);
  lbl4_g7924 : INR3D0BWP7T port map(A1 => lbl4_n_68, B1 => y_address(2), B2 => lbl4_n_21, ZN => lbl4_n_92);
  lbl4_g7926 : IND3D0BWP7T port map(A1 => lbl4_n_47, B1 => lbl4_n_31, B2 => lbl4_n_69, ZN => lbl4_n_86);
  lbl4_g7928 : AOI21D0BWP7T port map(A1 => lbl4_n_48, A2 => lbl4_n_12, B => lbl4_n_81, ZN => lbl4_n_89);
  lbl4_g7929 : OAI32D1BWP7T port map(A1 => lbl4_n_6, A2 => lbl4_n_32, A3 => lbl4_n_41, B1 => lbl4_n_26, B2 => lbl4_n_61, ZN => lbl4_n_88);
  lbl4_g7930 : AOI32D1BWP7T port map(A1 => lbl4_n_3, A2 => lbl4_n_42, A3 => lbl4_n_37, B1 => lbl4_n_69, B2 => lbl4_n_34, ZN => lbl4_n_87);
  lbl4_g7931 : OAI211D0BWP7T port map(A1 => lbl4_n_7, A2 => lbl4_n_19, B => lbl4_n_16, C => lbl4_n_35, ZN => lbl4_n_79);
  lbl4_g7932 : IND2D0BWP7T port map(A1 => lbl4_n_71, B1 => lbl4_n_6, ZN => lbl4_n_84);
  lbl4_g7933 : AOI21D0BWP7T port map(A1 => lbl4_n_53, A2 => x_address(1), B => lbl4_n_50, ZN => lbl4_n_83);
  lbl4_g7934 : NR2D0BWP7T port map(A1 => lbl4_n_27, A2 => lbl4_n_62, ZN => lbl4_n_82);
  lbl4_g7935 : IND2D1BWP7T port map(A1 => lbl4_n_52, B1 => lbl4_n_69, ZN => lbl4_n_81);
  lbl4_g7936 : IND2D1BWP7T port map(A1 => lbl4_n_48, B1 => lbl4_n_68, ZN => lbl4_n_80);
  lbl4_g7937 : OAI32D0BWP7T port map(A1 => x_address(2), A2 => lbl4_n_36, A3 => lbl4_n_19, B1 => x_address(1), B2 => lbl4_n_55, ZN => lbl4_n_73);
  lbl4_g7938 : IAO21D0BWP7T port map(A1 => lbl4_n_59, A2 => lbl4_n_8, B => y_address(4), ZN => lbl4_n_72);
  lbl4_g7939 : MOAI22D0BWP7T port map(A1 => lbl4_n_56, A2 => lbl4_n_18, B1 => lbl4_n_53, B2 => lbl4_n_13, ZN => lbl4_n_78);
  lbl4_g7940 : AOI32D1BWP7T port map(A1 => lbl4_n_31, A2 => y_address(2), A3 => y_address(1), B1 => lbl4_n_40, B2 => lbl4_n_25, ZN => lbl4_n_77);
  lbl4_g7941 : OA32D0BWP7T port map(A1 => y_address(3), A2 => lbl4_n_5, A3 => lbl4_n_23, B1 => lbl4_n_8, B2 => lbl4_n_41, Z => lbl4_n_76);
  lbl4_g7942 : AOI22D0BWP7T port map(A1 => lbl4_n_60, A2 => lbl4_n_13, B1 => lbl4_n_51, B2 => lbl4_n_19, ZN => lbl4_n_75);
  lbl4_g7943 : AO21D0BWP7T port map(A1 => lbl4_n_51, A2 => lbl4_n_9, B => lbl4_n_50, Z => lbl4_n_74);
  lbl4_g7944 : ND2D0BWP7T port map(A1 => lbl4_n_60, A2 => x_address(1), ZN => lbl4_n_67);
  lbl4_g7945 : ND2D0BWP7T port map(A1 => lbl4_n_40, A2 => lbl4_n_8, ZN => lbl4_n_71);
  lbl4_g7946 : NR2D0BWP7T port map(A1 => lbl4_n_58, A2 => x_address(1), ZN => lbl4_n_70);
  lbl4_g7947 : NR2D1BWP7T port map(A1 => map_selected(1), A2 => lbl4_n_56, ZN => lbl4_n_69);
  lbl4_g7948 : NR2D1BWP7T port map(A1 => lbl4_n_3, A2 => lbl4_n_52, ZN => lbl4_n_68);
  lbl4_g7949 : AOI32D0BWP7T port map(A1 => lbl4_n_5, A2 => lbl4_n_8, A3 => y_address(4), B1 => lbl4_n_16, B2 => y_address(3), ZN => lbl4_n_62);
  lbl4_g7950 : IND3D0BWP7T port map(A1 => lbl4_n_38, B1 => y_address(3), B2 => lbl4_n_11, ZN => lbl4_n_66);
  lbl4_g7951 : IAO21D0BWP7T port map(A1 => lbl4_n_30, A2 => lbl4_n_17, B => lbl4_n_53, ZN => lbl4_n_65);
  lbl4_g7952 : OR2D1BWP7T port map(A1 => lbl4_n_49, A2 => y_address(2), Z => lbl4_n_64);
  lbl4_g7953 : NR2D0BWP7T port map(A1 => lbl4_n_46, A2 => lbl4_n_15, ZN => lbl4_n_63);
  lbl4_g7954 : INVD0BWP7T port map(I => lbl4_n_58, ZN => lbl4_n_57);
  lbl4_g7956 : IND2D0BWP7T port map(A1 => lbl4_n_23, B1 => lbl4_n_16, ZN => lbl4_n_61);
  lbl4_g7957 : NR2D0BWP7T port map(A1 => lbl4_n_17, A2 => x_address(2), ZN => lbl4_n_60);
  lbl4_g7958 : IND2D0BWP7T port map(A1 => lbl4_n_29, B1 => y_address(2), ZN => lbl4_n_59);
  lbl4_g7959 : ND2D0BWP7T port map(A1 => lbl4_n_35, A2 => x_address(2), ZN => lbl4_n_58);
  lbl4_g7960 : IND2D0BWP7T port map(A1 => lbl4_n_17, B1 => x_address(2), ZN => lbl4_n_56);
  lbl4_g7961 : IND2D0BWP7T port map(A1 => lbl4_n_36, B1 => x_address(2), ZN => lbl4_n_55);
  lbl4_g7962 : INR2D0BWP7T port map(A1 => lbl4_n_30, B1 => lbl4_n_36, ZN => lbl4_n_54);
  lbl4_g7963 : INR2D0BWP7T port map(A1 => lbl4_n_37, B1 => x_address(2), ZN => lbl4_n_53);
  lbl4_g7964 : ND2D1BWP7T port map(A1 => lbl4_n_25, A2 => y_address(4), ZN => lbl4_n_52);
  lbl4_g7965 : INR2D0BWP7T port map(A1 => lbl4_n_37, B1 => lbl4_n_7, ZN => lbl4_n_51);
  lbl4_g7966 : INVD1BWP7T port map(I => lbl4_n_43, ZN => lbl4_n_42);
  lbl4_g7967 : INVD0BWP7T port map(I => lbl4_n_41, ZN => lbl4_n_40);
  lbl4_g7968 : ND2D1BWP7T port map(A1 => start_position_1(3), A2 => lbl4_n_27, ZN => start_position_0(2));
  lbl4_g7969 : INR2D0BWP7T port map(A1 => lbl4_n_30, B1 => lbl4_n_17, ZN => lbl4_n_50);
  lbl4_g7970 : OR2D1BWP7T port map(A1 => lbl4_n_22, A2 => lbl4_n_26, Z => lbl4_n_49);
  lbl4_g7971 : MAOI22D0BWP7T port map(A1 => lbl4_n_5, A2 => y_address(1), B1 => lbl4_n_5, B2 => y_address(1), ZN => lbl4_n_48);
  lbl4_g7972 : INR2D0BWP7T port map(A1 => lbl4_n_20, B1 => lbl4_n_13, ZN => lbl4_n_47);
  lbl4_g7973 : INR2D0BWP7T port map(A1 => lbl4_n_21, B1 => lbl4_n_11, ZN => lbl4_n_46);
  lbl4_g7974 : ND2D0BWP7T port map(A1 => lbl4_n_30, A2 => lbl4_n_37, ZN => lbl4_n_45);
  lbl4_g7975 : NR3D0BWP7T port map(A1 => lbl4_n_7, A2 => lbl4_n_9, A3 => x_address(3), ZN => lbl4_n_44);
  lbl4_g7976 : ND2D0BWP7T port map(A1 => lbl4_n_30, A2 => lbl4_n_4, ZN => lbl4_n_43);
  lbl4_g7977 : ND2D0BWP7T port map(A1 => lbl4_n_29, A2 => lbl4_n_5, ZN => lbl4_n_41);
  lbl4_g7978 : CKND1BWP7T port map(I => lbl4_n_34, ZN => lbl4_n_33);
  lbl4_g7979 : INVD1BWP7T port map(I => lbl4_n_32, ZN => lbl4_n_31);
  lbl4_g7980 : INVD1BWP7T port map(I => start_position_0(3), ZN => lbl4_n_27);
  lbl4_g7981 : INVD1BWP7T port map(I => lbl4_n_26, ZN => lbl4_n_25);
  lbl4_g7982 : ND2D0BWP7T port map(A1 => y_address(2), A2 => y_address(4), ZN => lbl4_n_38);
  lbl4_g7983 : INR2D0BWP7T port map(A1 => x_address(4), B1 => x_address(3), ZN => lbl4_n_37);
  lbl4_g7984 : ND2D0BWP7T port map(A1 => x_address(3), A2 => x_address(4), ZN => lbl4_n_36);
  lbl4_g7985 : NR2D0BWP7T port map(A1 => x_address(4), A2 => x_address(3), ZN => lbl4_n_35);
  lbl4_g7986 : NR2D0BWP7T port map(A1 => lbl4_n_4, A2 => lbl4_n_9, ZN => lbl4_n_34);
  lbl4_g7987 : ND2D1BWP7T port map(A1 => map_selected(0), A2 => lbl4_n_8, ZN => lbl4_n_32);
  lbl4_g7988 : NR2D0BWP7T port map(A1 => x_address(2), A2 => x_address(1), ZN => lbl4_n_30);
  lbl4_g7989 : NR2D0BWP7T port map(A1 => y_address(1), A2 => y_address(0), ZN => lbl4_n_29);
  lbl4_g7990 : NR2D1BWP7T port map(A1 => lbl4_n_3, A2 => map_selected(0), ZN => start_position_0(3));
  lbl4_g7991 : ND2D1BWP7T port map(A1 => map_selected(0), A2 => y_address(3), ZN => lbl4_n_26);
  lbl4_g7992 : INVD0BWP7T port map(I => lbl4_n_18, ZN => lbl4_n_19);
  lbl4_g7993 : INVD1BWP7T port map(I => lbl4_n_16, ZN => lbl4_n_15);
  lbl4_g7994 : INVD1BWP7T port map(I => lbl4_n_14, ZN => lbl4_n_13);
  lbl4_g7995 : INVD1BWP7T port map(I => lbl4_n_12, ZN => lbl4_n_11);
  lbl4_g7996 : ND2D0BWP7T port map(A1 => map_selected(1), A2 => map_selected(0), ZN => start_position_1(5));
  lbl4_g7997 : ND2D1BWP7T port map(A1 => lbl4_n_3, A2 => map_selected(0), ZN => start_position_1(3));
  lbl4_g7998 : ND2D0BWP7T port map(A1 => y_address(1), A2 => y_address(0), ZN => lbl4_n_23);
  lbl4_g7999 : ND2D1BWP7T port map(A1 => map_selected(1), A2 => lbl4_n_6, ZN => lbl4_n_22);
  lbl4_g8000 : IND2D0BWP7T port map(A1 => y_address(0), B1 => y_address(1), ZN => lbl4_n_21);
  lbl4_g8001 : ND2D0BWP7T port map(A1 => lbl4_n_9, A2 => x_address(0), ZN => lbl4_n_20);
  lbl4_g8002 : ND2D0BWP7T port map(A1 => lbl4_n_4, A2 => lbl4_n_9, ZN => lbl4_n_18);
  lbl4_g8003 : IND2D0BWP7T port map(A1 => x_address(4), B1 => x_address(3), ZN => lbl4_n_17);
  lbl4_g8004 : NR2D0BWP7T port map(A1 => lbl4_n_5, A2 => y_address(4), ZN => lbl4_n_16);
  lbl4_g8005 : ND2D0BWP7T port map(A1 => lbl4_n_4, A2 => x_address(1), ZN => lbl4_n_14);
  lbl4_g8006 : IND2D0BWP7T port map(A1 => y_address(1), B1 => y_address(0), ZN => lbl4_n_12);
  lbl4_g8007 : INVD1BWP7T port map(I => x_address(1), ZN => lbl4_n_9);
  lbl4_g8008 : INVD1BWP7T port map(I => y_address(3), ZN => lbl4_n_8);
  lbl4_g8009 : INVD0BWP7T port map(I => x_address(2), ZN => lbl4_n_7);
  lbl4_g8010 : INVD1BWP7T port map(I => y_address(4), ZN => lbl4_n_6);
  lbl4_g8011 : INVD1BWP7T port map(I => y_address(2), ZN => lbl4_n_5);
  lbl4_g8012 : INVD1BWP7T port map(I => x_address(0), ZN => lbl4_n_4);
  lbl4_g8013 : INVD1BWP7T port map(I => map_selected(1), ZN => lbl4_n_3);
  lbl4_g8014 : AO32D1BWP7T port map(A1 => lbl4_n_70, A2 => lbl4_n_63, A3 => lbl4_n_25, B1 => lbl4_n_88, B2 => lbl4_n_54, Z => lbl4_n_161);
  lbl2_dec1_g100 : AO22D0BWP7T port map(A1 => lbl2_dec1_n_2, A2 => lbl2_data_synced(4), B1 => lbl2_data_synced(5), B2 => lbl2_dec1_n_1, Z => lbl2_walls(6));
  lbl2_dec1_g101 : IOA21D1BWP7T port map(A1 => lbl2_dec1_n_2, A2 => lbl2_dec1_n_0, B => lbl2_dec1_n_5, ZN => lbl2_walls(4));
  lbl2_dec1_g102 : IND2D1BWP7T port map(A1 => lbl2_dec1_n_2, B1 => lbl2_dec1_n_3, ZN => lbl2_walls(5));
  lbl2_dec1_g103 : IOA21D1BWP7T port map(A1 => lbl2_dec1_n_0, A2 => lbl2_data_synced(6), B => lbl2_data_synced(5), ZN => lbl2_dec1_n_5);
  lbl2_dec1_g104 : IOA21D1BWP7T port map(A1 => lbl2_data_synced(6), A2 => lbl2_data_synced(5), B => lbl2_dec1_n_3, ZN => lbl2_walls(7));
  lbl2_dec1_g105 : IND2D1BWP7T port map(A1 => lbl2_data_synced(6), B1 => lbl2_data_synced(4), ZN => lbl2_dec1_n_3);
  lbl2_dec1_g106 : ND2D0BWP7T port map(A1 => lbl2_data_synced(6), A2 => lbl2_data_synced(4), ZN => lbl2_dec1_n_1);
  lbl2_dec1_g107 : INR2D1BWP7T port map(A1 => lbl2_data_synced(6), B1 => lbl2_data_synced(5), ZN => lbl2_dec1_n_2);
  lbl2_dec1_g108 : INVD0BWP7T port map(I => lbl2_data_synced(4), ZN => lbl2_dec1_n_0);
  lbl2_hscr_g18635 : IOA21D1BWP7T port map(A1 => lbl2_pixelator_color(3), A2 => lbl2_hscr_n_203, B => lbl2_hscr_n_370, ZN => lbl2_homescreen_color(3));
  lbl2_hscr_g18636 : IOA21D1BWP7T port map(A1 => lbl2_pixelator_color(2), A2 => lbl2_hscr_n_203, B => lbl2_hscr_n_370, ZN => lbl2_homescreen_color(2));
  lbl2_hscr_g18637 : IOA21D1BWP7T port map(A1 => lbl2_pixelator_color(1), A2 => lbl2_hscr_n_203, B => lbl2_hscr_n_371, ZN => lbl2_homescreen_color(1));
  lbl2_hscr_g18638 : IOA21D1BWP7T port map(A1 => lbl2_pixelator_color(0), A2 => lbl2_hscr_n_203, B => lbl2_hscr_n_371, ZN => lbl2_homescreen_color(0));
  lbl2_hscr_g18639 : IOA21D1BWP7T port map(A1 => lbl2_hscr_n_368, A2 => lbl2_hscr_n_345, B => lbl2_hscr_n_369, ZN => lbl2_hscr_n_371);
  lbl2_hscr_g18640 : IOA21D1BWP7T port map(A1 => lbl2_hscr_n_368, A2 => lbl2_hscr_n_328, B => lbl2_hscr_n_369, ZN => lbl2_hscr_n_370);
  lbl2_hscr_g18641 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_368, A2 => lbl2_hscr_n_360, B => lbl2_hscr_n_203, ZN => lbl2_hscr_n_369);
  lbl2_hscr_g18642 : AOI222D0BWP7T port map(A1 => lbl2_hscr_n_367, A2 => lbl2_hscr_n_180, B1 => lbl2_hscr_n_348, B2 => lbl2_hscr_n_32, C1 => lbl2_hscr_n_247, C2 => lbl2_hscr_n_110, ZN => lbl2_hscr_n_368);
  lbl2_hscr_g18643 : AOI211D1BWP7T port map(A1 => lbl2_hscr_n_10, A2 => lbl2_v_count(4), B => lbl2_hscr_n_366, C => lbl2_hscr_n_59, ZN => lbl2_hscr_n_367);
  lbl2_hscr_g18644 : OAI211D1BWP7T port map(A1 => lbl2_v_count(5), A2 => lbl2_hscr_n_10, B => lbl2_hscr_n_365, C => lbl2_hscr_n_38, ZN => lbl2_hscr_n_366);
  lbl2_hscr_g18645 : AO211D0BWP7T port map(A1 => lbl2_hscr_n_191, A2 => lbl2_hscr_n_198, B => lbl2_hscr_n_364, C => lbl2_hscr_n_291, Z => lbl2_hscr_n_365);
  lbl2_hscr_g18646 : IND4D0BWP7T port map(A1 => lbl2_hscr_n_363, B1 => lbl2_hscr_n_266, B2 => lbl2_hscr_n_344, B3 => lbl2_hscr_n_355, ZN => lbl2_hscr_n_364);
  lbl2_hscr_g18647 : ND4D0BWP7T port map(A1 => lbl2_hscr_n_362, A2 => lbl2_hscr_n_359, A3 => lbl2_hscr_n_361, A4 => lbl2_hscr_n_358, ZN => lbl2_hscr_n_363);
  lbl2_hscr_g18648 : OAI31D0BWP7T port map(A1 => lbl2_hscr_n_256, A2 => lbl2_hscr_n_321, A3 => lbl2_hscr_n_357, B => lbl2_h_count(0), ZN => lbl2_hscr_n_362);
  lbl2_hscr_g18649 : OAI31D0BWP7T port map(A1 => lbl2_hscr_n_210, A2 => lbl2_hscr_n_299, A3 => lbl2_hscr_n_350, B => FE_DBTN1_lbl2_h_count_1, ZN => lbl2_hscr_n_361);
  lbl2_hscr_g18650 : ND4D0BWP7T port map(A1 => lbl2_hscr_n_349, A2 => lbl2_hscr_n_73, A3 => lbl2_hscr_n_35, A4 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_360);
  lbl2_hscr_g18651 : NR4D0BWP7T port map(A1 => lbl2_hscr_n_352, A2 => lbl2_hscr_n_356, A3 => lbl2_hscr_n_343, A4 => lbl2_hscr_n_325, ZN => lbl2_hscr_n_359);
  lbl2_hscr_g18652 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_306, A2 => lbl2_hscr_n_103, B1 => lbl2_hscr_n_239, B2 => lbl2_hscr_n_71, C => lbl2_hscr_n_354, ZN => lbl2_hscr_n_358);
  lbl2_hscr_g18653 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_143, A2 => lbl2_hscr_n_209, B => lbl2_hscr_n_353, C => lbl2_hscr_n_212, ZN => lbl2_hscr_n_357);
  lbl2_hscr_g18654 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_351, A2 => FE_DBTN1_lbl2_h_count_1, ZN => lbl2_hscr_n_356);
  lbl2_hscr_g18655 : OAI31D0BWP7T port map(A1 => lbl2_hscr_n_257, A2 => lbl2_hscr_n_290, A3 => lbl2_hscr_n_341, B => lbl2_h_count(2), ZN => lbl2_hscr_n_355);
  lbl2_hscr_g18656 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_347, A2 => lbl2_h_count(2), B1 => lbl2_hscr_n_208, B2 => lbl2_hscr_n_138, ZN => lbl2_hscr_n_354);
  lbl2_hscr_g18657 : MAOI22D0BWP7T port map(A1 => lbl2_hscr_n_288, A2 => lbl2_hscr_n_103, B1 => lbl2_hscr_n_346, B2 => FE_DBTN1_lbl2_h_count_1, ZN => lbl2_hscr_n_353);
  lbl2_hscr_g18658 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_333, A2 => lbl2_hscr_n_300, A3 => lbl2_hscr_n_223, B => lbl2_h_count(0), ZN => lbl2_hscr_n_352);
  lbl2_hscr_g18659 : NR4D0BWP7T port map(A1 => lbl2_hscr_n_336, A2 => lbl2_hscr_n_321, A3 => lbl2_hscr_n_282, A4 => lbl2_hscr_n_256, ZN => lbl2_hscr_n_351);
  lbl2_hscr_g18660 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_82, A2 => lbl2_hscr_n_242, B => lbl2_hscr_n_342, C => lbl2_hscr_n_223, ZN => lbl2_hscr_n_350);
  lbl2_hscr_g18661 : MAOI22D0BWP7T port map(A1 => lbl2_hscr_n_51, A2 => lbl2_v_count(6), B1 => lbl2_hscr_n_345, B2 => lbl2_hscr_n_328, ZN => lbl2_hscr_n_349);
  lbl2_hscr_g18662 : AOI211D1BWP7T port map(A1 => lbl2_hscr_n_308, A2 => lbl2_hscr_n_6, B => lbl2_hscr_n_338, C => lbl2_hscr_n_58, ZN => lbl2_hscr_n_348);
  lbl2_hscr_g18663 : NR4D0BWP7T port map(A1 => lbl2_hscr_n_330, A2 => lbl2_hscr_n_302, A3 => lbl2_hscr_n_292, A4 => lbl2_hscr_n_270, ZN => lbl2_hscr_n_347);
  lbl2_hscr_g18664 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_273, A2 => lbl2_hscr_n_3, B1 => lbl2_hscr_n_293, B2 => lbl2_hscr_n_156, C => lbl2_hscr_n_339, ZN => lbl2_hscr_n_346);
  lbl2_hscr_g18665 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_269, A2 => lbl2_hscr_n_116, B1 => lbl2_hscr_n_253, B2 => lbl2_v_count(1), C => lbl2_hscr_n_334, ZN => lbl2_hscr_n_344);
  lbl2_hscr_g18666 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_161, A2 => lbl2_hscr_n_244, B => lbl2_hscr_n_335, C => lbl2_hscr_n_276, ZN => lbl2_hscr_n_345);
  lbl2_hscr_g18667 : OA31D1BWP7T port map(A1 => lbl2_hscr_n_257, A2 => lbl2_hscr_n_283, A3 => lbl2_hscr_n_326, B => lbl2_hscr_n_29, Z => lbl2_hscr_n_343);
  lbl2_hscr_g18668 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_250, A2 => lbl2_hscr_n_120, B1 => lbl2_hscr_n_232, B2 => lbl2_hscr_n_133, C => lbl2_hscr_n_340, ZN => lbl2_hscr_n_342);
  lbl2_hscr_g18669 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_206, A2 => lbl2_hscr_n_47, B => lbl2_hscr_n_337, ZN => lbl2_hscr_n_341);
  lbl2_hscr_g18670 : OAI211D1BWP7T port map(A1 => lbl2_v_count(0), A2 => lbl2_hscr_n_233, B => lbl2_hscr_n_327, C => lbl2_hscr_n_296, ZN => lbl2_hscr_n_340);
  lbl2_hscr_g18671 : ND4D0BWP7T port map(A1 => lbl2_hscr_n_322, A2 => lbl2_hscr_n_286, A3 => lbl2_hscr_n_261, A4 => lbl2_hscr_n_260, ZN => lbl2_hscr_n_339);
  lbl2_hscr_g18672 : IND4D0BWP7T port map(A1 => lbl2_v_count(5), B1 => lbl2_v_count(8), B2 => lbl2_hscr_n_26, B3 => lbl2_hscr_n_320, ZN => lbl2_hscr_n_338);
  lbl2_hscr_g18673 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_317, A2 => lbl2_hscr_n_47, B1 => lbl2_hscr_n_168, B2 => lbl2_hscr_n_183, C => lbl2_hscr_n_210, ZN => lbl2_hscr_n_337);
  lbl2_hscr_g18674 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_123, A2 => lbl2_hscr_n_274, B => lbl2_hscr_n_323, C => lbl2_hscr_n_304, ZN => lbl2_hscr_n_336);
  lbl2_hscr_g18675 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_204, A2 => lbl2_hscr_n_198, A3 => lbl2_hscr_n_25, B => lbl2_hscr_n_331, ZN => lbl2_hscr_n_335);
  lbl2_hscr_g18676 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_226, A2 => lbl2_hscr_n_147, B => lbl2_hscr_n_329, C => lbl2_hscr_n_215, ZN => lbl2_hscr_n_334);
  lbl2_hscr_g18677 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_210, A2 => lbl2_v_count(0), B => lbl2_hscr_n_332, ZN => lbl2_hscr_n_333);
  lbl2_hscr_g18678 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_164, A2 => lbl2_hscr_n_200, B => lbl2_hscr_n_324, C => lbl2_hscr_n_211, ZN => lbl2_hscr_n_332);
  lbl2_hscr_g18679 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_315, A2 => lbl2_hscr_n_48, B => lbl2_hscr_n_316, ZN => lbl2_hscr_n_331);
  lbl2_hscr_g18680 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_298, A2 => lbl2_hscr_n_259, A3 => lbl2_hscr_n_255, B => lbl2_hscr_n_47, ZN => lbl2_hscr_n_330);
  lbl2_hscr_g18681 : AOI211XD0BWP7T port map(A1 => lbl2_hscr_n_163, A2 => lbl2_hscr_n_182, B => lbl2_hscr_n_313, C => lbl2_hscr_n_301, ZN => lbl2_hscr_n_329);
  lbl2_hscr_g18682 : OA221D0BWP7T port map(A1 => lbl2_hscr_n_207, A2 => lbl2_hscr_n_158, B1 => lbl2_hscr_n_142, B2 => lbl2_hscr_n_208, C => lbl2_hscr_n_314, Z => lbl2_hscr_n_327);
  lbl2_hscr_g18683 : OAI31D0BWP7T port map(A1 => lbl2_hscr_n_68, A2 => lbl2_hscr_n_145, A3 => lbl2_hscr_n_243, B => lbl2_hscr_n_319, ZN => lbl2_hscr_n_326);
  lbl2_hscr_g18684 : OAI221D0BWP7T port map(A1 => lbl2_hscr_n_271, A2 => lbl2_hscr_n_145, B1 => lbl2_hscr_n_91, B2 => lbl2_hscr_n_246, C => lbl2_hscr_n_318, ZN => lbl2_hscr_n_328);
  lbl2_hscr_g18685 : AOI211D1BWP7T port map(A1 => lbl2_hscr_n_305, A2 => lbl2_hscr_n_233, B => lbl2_h_count(1), C => lbl2_hscr_n_9, ZN => lbl2_hscr_n_325);
  lbl2_hscr_g18686 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_234, A2 => lbl2_hscr_n_103, A3 => lbl2_hscr_n_47, B1 => lbl2_hscr_n_309, B2 => lbl2_h_count(1), ZN => lbl2_hscr_n_324);
  lbl2_hscr_g18687 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_175, A2 => lbl2_hscr_n_116, A3 => lbl2_hscr_n_71, B1 => lbl2_hscr_n_310, B2 => lbl2_hscr_n_103, ZN => lbl2_hscr_n_323);
  lbl2_hscr_g18688 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_303, A2 => lbl2_h_count(2), B1 => lbl2_hscr_n_251, B2 => lbl2_hscr_n_122, ZN => lbl2_hscr_n_322);
  lbl2_hscr_g18689 : AOI211D1BWP7T port map(A1 => lbl2_v_count(2), A2 => lbl2_v_count(4), B => lbl2_hscr_n_311, C => lbl2_hscr_n_238, ZN => lbl2_hscr_n_320);
  lbl2_hscr_g18690 : OA221D0BWP7T port map(A1 => lbl2_hscr_n_200, A2 => lbl2_hscr_n_141, B1 => lbl2_hscr_n_121, B2 => lbl2_hscr_n_208, C => lbl2_hscr_n_307, Z => lbl2_hscr_n_319);
  lbl2_hscr_g18691 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_236, A2 => lbl2_hscr_n_192, B1 => lbl2_hscr_n_267, B2 => lbl2_hscr_n_159, C => lbl2_hscr_n_294, ZN => lbl2_hscr_n_318);
  lbl2_hscr_g18692 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_155, A2 => lbl2_hscr_n_184, B => lbl2_hscr_n_280, C => lbl2_hscr_n_264, ZN => lbl2_hscr_n_321);
  lbl2_hscr_g18693 : AO221D0BWP7T port map(A1 => lbl2_hscr_n_195, A2 => lbl2_hscr_n_159, B1 => lbl2_hscr_n_269, B2 => lbl2_hscr_n_64, C => lbl2_hscr_n_187, Z => lbl2_hscr_n_317);
  lbl2_hscr_g18694 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_275, A2 => lbl2_hscr_n_159, A3 => lbl2_hscr_n_48, B1 => lbl2_hscr_n_284, B2 => lbl2_hscr_n_180, ZN => lbl2_hscr_n_316);
  lbl2_hscr_g18695 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_221, A2 => lbl2_hscr_n_114, A3 => lbl2_hscr_n_116, B => lbl2_hscr_n_312, ZN => lbl2_hscr_n_315);
  lbl2_hscr_g18696 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_289, A2 => lbl2_hscr_n_71, B1 => lbl2_hscr_n_199, B2 => lbl2_hscr_n_169, ZN => lbl2_hscr_n_314);
  lbl2_hscr_g18697 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_295, A2 => lbl2_hscr_n_90, B1 => lbl2_hscr_n_262, B2 => lbl2_hscr_n_47, ZN => lbl2_hscr_n_313);
  lbl2_hscr_g18698 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_244, A2 => lbl2_hscr_n_64, B => lbl2_hscr_n_285, ZN => lbl2_hscr_n_312);
  lbl2_hscr_g18699 : OAI31D0BWP7T port map(A1 => direction_in(3), A2 => lbl2_hscr_n_66, A3 => lbl2_hscr_n_278, B => lbl2_hscr_n_150, ZN => lbl2_hscr_n_311);
  lbl2_hscr_g18700 : AO211D0BWP7T port map(A1 => lbl2_hscr_n_227, A2 => lbl2_hscr_n_98, B => lbl2_hscr_n_288, C => lbl2_hscr_n_224, Z => lbl2_hscr_n_310);
  lbl2_hscr_g18701 : OAI221D0BWP7T port map(A1 => lbl2_hscr_n_233, A2 => lbl2_hscr_n_2, B1 => lbl2_hscr_n_47, B2 => lbl2_hscr_n_255, C => lbl2_hscr_n_287, ZN => lbl2_hscr_n_309);
  lbl2_hscr_g18702 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_278, A2 => direction_in(2), B => lbl2_central_x_vec(8), ZN => lbl2_hscr_n_308);
  lbl2_hscr_g18703 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_194, A2 => lbl2_hscr_n_118, A3 => lbl2_hscr_n_71, B => lbl2_hscr_n_281, ZN => lbl2_hscr_n_307);
  lbl2_hscr_g18704 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_117, A2 => lbl2_hscr_n_229, B => lbl2_hscr_n_245, C => lbl2_hscr_n_265, ZN => lbl2_hscr_n_306);
  lbl2_hscr_g18705 : AOI222D0BWP7T port map(A1 => lbl2_hscr_n_199, A2 => lbl2_hscr_n_140, B1 => lbl2_hscr_n_250, B2 => lbl2_hscr_n_97, C1 => lbl2_hscr_n_254, C2 => lbl2_hscr_n_64, ZN => lbl2_hscr_n_305);
  lbl2_hscr_g18706 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_263, A2 => lbl2_hscr_n_3, B1 => lbl2_hscr_n_199, B2 => lbl2_hscr_n_178, ZN => lbl2_hscr_n_304);
  lbl2_hscr_g18707 : AO21D0BWP7T port map(A1 => lbl2_hscr_n_182, A2 => lbl2_hscr_n_137, B => lbl2_hscr_n_297, Z => lbl2_hscr_n_303);
  lbl2_hscr_g18708 : OAI32D1BWP7T port map(A1 => lbl2_hscr_n_101, A2 => lbl2_hscr_n_134, A3 => lbl2_hscr_n_193, B1 => lbl2_hscr_n_96, B2 => lbl2_hscr_n_279, ZN => lbl2_hscr_n_302);
  lbl2_hscr_g18709 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_279, A2 => lbl2_hscr_n_124, B1 => lbl2_hscr_n_214, B2 => lbl2_v_count(1), ZN => lbl2_hscr_n_301);
  lbl2_hscr_g18710 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_277, A2 => lbl2_hscr_n_47, B1 => lbl2_hscr_n_250, B2 => lbl2_hscr_n_176, ZN => lbl2_hscr_n_300);
  lbl2_hscr_g18711 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_268, A2 => lbl2_hscr_n_91, B1 => lbl2_hscr_n_220, B2 => lbl2_hscr_n_48, ZN => lbl2_hscr_n_299);
  lbl2_hscr_g18712 : OA22D0BWP7T port map(A1 => lbl2_hscr_n_272, A2 => lbl2_hscr_n_161, B1 => lbl2_hscr_n_138, B2 => lbl2_hscr_n_226, Z => lbl2_hscr_n_298);
  lbl2_hscr_g18713 : AOI211D1BWP7T port map(A1 => lbl2_hscr_n_228, A2 => lbl2_hscr_n_229, B => lbl2_hscr_n_117, C => lbl2_hscr_n_82, ZN => lbl2_hscr_n_297);
  lbl2_hscr_g18714 : IND4D0BWP7T port map(A1 => lbl2_hscr_n_124, B1 => lbl2_h_count(2), B2 => lbl2_v_count(1), B3 => lbl2_hscr_n_227, ZN => lbl2_hscr_n_296);
  lbl2_hscr_g18715 : OA211D0BWP7T port map(A1 => lbl2_hscr_n_99, A2 => lbl2_hscr_n_226, B => lbl2_hscr_n_245, C => lbl2_hscr_n_222, Z => lbl2_hscr_n_295);
  lbl2_hscr_g18716 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_246, A2 => lbl2_hscr_n_116, A3 => lbl2_hscr_n_82, ZN => lbl2_hscr_n_294);
  lbl2_hscr_g18717 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_243, A2 => lbl2_hscr_n_83, B => lbl2_hscr_n_173, ZN => lbl2_hscr_n_293);
  lbl2_hscr_g18718 : AOI211D1BWP7T port map(A1 => lbl2_hscr_n_243, A2 => lbl2_hscr_n_173, B => lbl2_hscr_n_101, C => lbl2_hscr_n_145, ZN => lbl2_hscr_n_292);
  lbl2_hscr_g18719 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_242, A2 => lbl2_hscr_n_235, B => lbl2_hscr_n_91, ZN => lbl2_hscr_n_291);
  lbl2_hscr_g18720 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_242, A2 => lbl2_hscr_n_82, A3 => lbl2_hscr_n_83, ZN => lbl2_hscr_n_290);
  lbl2_hscr_g18721 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_234, B1 => lbl2_hscr_n_258, ZN => lbl2_hscr_n_289);
  lbl2_hscr_g18722 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_250, A2 => lbl2_hscr_n_140, B1 => lbl2_hscr_n_199, B2 => lbl2_hscr_n_97, ZN => lbl2_hscr_n_287);
  lbl2_hscr_g18723 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_225, A2 => lbl2_hscr_n_153, A3 => lbl2_hscr_n_67, B1 => lbl2_hscr_n_232, B2 => lbl2_hscr_n_144, ZN => lbl2_hscr_n_286);
  lbl2_hscr_g18724 : AOI33D1BWP7T port map(A1 => lbl2_hscr_n_204, A2 => lbl2_hscr_n_216, A3 => lbl2_hscr_n_145, B1 => lbl2_hscr_n_194, B2 => lbl2_hscr_n_180, B3 => lbl2_hscr_n_51, ZN => lbl2_hscr_n_285);
  lbl2_hscr_g18725 : OAI33D1BWP7T port map(A1 => lbl2_hscr_n_47, A2 => lbl2_hscr_n_116, A3 => lbl2_hscr_n_218, B1 => lbl2_hscr_n_52, B2 => lbl2_hscr_n_171, B3 => lbl2_hscr_n_155, ZN => lbl2_hscr_n_284);
  lbl2_hscr_g18726 : OAI33D1BWP7T port map(A1 => lbl2_hscr_n_1, A2 => lbl2_hscr_n_82, A3 => lbl2_hscr_n_213, B1 => lbl2_hscr_n_3, B2 => lbl2_hscr_n_119, B3 => lbl2_hscr_n_229, ZN => lbl2_hscr_n_283);
  lbl2_hscr_g18727 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_209, A2 => lbl2_hscr_n_127, B1 => lbl2_hscr_n_249, B2 => lbl2_hscr_n_158, ZN => lbl2_hscr_n_282);
  lbl2_hscr_g18728 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_240, A2 => lbl2_hscr_n_230, B1 => lbl2_hscr_n_207, B2 => lbl2_hscr_n_148, ZN => lbl2_hscr_n_281);
  lbl2_hscr_g18729 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_250, A2 => lbl2_hscr_n_167, B1 => lbl2_hscr_n_232, B2 => lbl2_hscr_n_157, ZN => lbl2_hscr_n_280);
  lbl2_hscr_g18730 : OAI31D0BWP7T port map(A1 => lbl2_hscr_n_116, A2 => lbl2_hscr_n_135, A3 => lbl2_hscr_n_231, B => lbl2_hscr_n_235, ZN => lbl2_hscr_n_288);
  lbl2_hscr_g18731 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_230, A2 => lbl2_hscr_n_149, B => lbl2_hscr_n_220, ZN => lbl2_hscr_n_277);
  lbl2_hscr_g18732 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_230, B1 => lbl2_hscr_n_50, B2 => lbl2_hscr_n_180, ZN => lbl2_hscr_n_276);
  lbl2_hscr_g18733 : IOA21D1BWP7T port map(A1 => lbl2_hscr_n_221, A2 => lbl2_hscr_n_108, B => lbl2_hscr_n_217, ZN => lbl2_hscr_n_275);
  lbl2_hscr_g18734 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_183, A2 => lbl2_hscr_n_2, A3 => lbl2_h_count(2), B => lbl2_hscr_n_251, ZN => lbl2_hscr_n_274);
  lbl2_hscr_g18735 : OAI31D0BWP7T port map(A1 => lbl2_v_count(0), A2 => lbl2_hscr_n_101, A3 => lbl2_hscr_n_197, B => lbl2_hscr_n_252, ZN => lbl2_hscr_n_273);
  lbl2_hscr_g18736 : OA21D0BWP7T port map(A1 => lbl2_hscr_n_231, A2 => lbl2_hscr_n_104, B => lbl2_hscr_n_184, Z => lbl2_hscr_n_272);
  lbl2_hscr_g18737 : IND4D0BWP7T port map(A1 => lbl2_hscr_n_90, B1 => lbl2_hscr_n_76, B2 => lbl2_hscr_n_172, B3 => lbl2_hscr_n_205, ZN => lbl2_hscr_n_271);
  lbl2_hscr_g18738 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_228, A2 => lbl2_hscr_n_117, A3 => lbl2_hscr_n_1, ZN => lbl2_hscr_n_270);
  lbl2_hscr_g18739 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_226, A2 => lbl2_hscr_n_1, B => lbl2_hscr_n_202, ZN => lbl2_hscr_n_279);
  lbl2_hscr_g18740 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_9, A2 => lbl2_hscr_n_84, B => lbl2_hscr_n_248, C => lbl2_hscr_n_81, ZN => lbl2_hscr_n_278);
  lbl2_hscr_g18741 : INVD0BWP7T port map(I => lbl2_hscr_n_269, ZN => lbl2_hscr_n_268);
  lbl2_hscr_g18742 : AO22D0BWP7T port map(A1 => lbl2_hscr_n_236, A2 => lbl2_hscr_n_50, B1 => lbl2_hscr_n_108, B2 => lbl2_hscr_n_205, Z => lbl2_hscr_n_267);
  lbl2_hscr_g18743 : IOA21D1BWP7T port map(A1 => lbl2_hscr_n_138, A2 => lbl2_hscr_n_96, B => lbl2_hscr_n_251, ZN => lbl2_hscr_n_266);
  lbl2_hscr_g18744 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_231, A2 => lbl2_hscr_n_143, B => lbl2_hscr_n_241, ZN => lbl2_hscr_n_265);
  lbl2_hscr_g18745 : OA33D0BWP7T port map(A1 => lbl2_hscr_n_101, A2 => lbl2_hscr_n_172, A3 => lbl2_hscr_n_173, B1 => lbl2_v_count(1), B2 => lbl2_hscr_n_96, B3 => lbl2_hscr_n_201, Z => lbl2_hscr_n_264);
  lbl2_hscr_g18746 : OAI32D1BWP7T port map(A1 => lbl2_hscr_n_47, A2 => lbl2_hscr_n_134, A3 => lbl2_hscr_n_181, B1 => lbl2_hscr_n_124, B2 => lbl2_hscr_n_226, ZN => lbl2_hscr_n_263);
  lbl2_hscr_g18747 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_202, A2 => lbl2_hscr_n_137, B => lbl2_hscr_n_253, ZN => lbl2_hscr_n_262);
  lbl2_hscr_g18748 : OA22D0BWP7T port map(A1 => lbl2_hscr_n_237, A2 => lbl2_hscr_n_90, B1 => lbl2_hscr_n_48, B2 => lbl2_hscr_n_206, Z => lbl2_hscr_n_261);
  lbl2_hscr_g18749 : OA22D0BWP7T port map(A1 => lbl2_hscr_n_222, A2 => lbl2_hscr_n_102, B1 => lbl2_hscr_n_96, B2 => lbl2_hscr_n_209, Z => lbl2_hscr_n_260);
  lbl2_hscr_g18750 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_0, A2 => lbl2_hscr_n_82, B1 => lbl2_hscr_n_202, B2 => lbl2_hscr_n_122, ZN => lbl2_hscr_n_259);
  lbl2_hscr_g18751 : MAOI22D0BWP7T port map(A1 => lbl2_hscr_n_227, A2 => lbl2_hscr_n_118, B1 => lbl2_hscr_n_154, B2 => lbl2_hscr_n_142, ZN => lbl2_hscr_n_258);
  lbl2_hscr_g18752 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_193, A2 => lbl2_hscr_n_125, B1 => lbl2_hscr_n_229, B2 => lbl2_hscr_n_106, ZN => lbl2_hscr_n_269);
  lbl2_hscr_g18753 : INVD0BWP7T port map(I => lbl2_hscr_n_255, ZN => lbl2_hscr_n_254);
  lbl2_hscr_g18754 : INVD0BWP7T port map(I => lbl2_hscr_n_252, ZN => lbl2_hscr_n_253);
  lbl2_hscr_g18755 : INVD0BWP7T port map(I => lbl2_hscr_n_250, ZN => lbl2_hscr_n_249);
  lbl2_hscr_g18756 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_126, A2 => lbl2_h_count(2), B => lbl2_hscr_n_219, ZN => lbl2_hscr_n_248);
  lbl2_hscr_g18757 : OAI31D0BWP7T port map(A1 => lbl2_h_count(4), A2 => lbl2_h_count(2), A3 => lbl2_hscr_n_177, B => lbl2_hscr_n_185, ZN => lbl2_hscr_n_247);
  lbl2_hscr_g18758 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_170, A2 => lbl2_hscr_n_228, ZN => lbl2_hscr_n_257);
  lbl2_hscr_g18759 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_190, A2 => lbl2_hscr_n_47, A3 => lbl2_h_count(2), ZN => lbl2_hscr_n_256);
  lbl2_hscr_g18760 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_231, B1 => lbl2_hscr_n_137, ZN => lbl2_hscr_n_255);
  lbl2_hscr_g18761 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_226, B1 => lbl2_hscr_n_118, ZN => lbl2_hscr_n_252);
  lbl2_hscr_g18762 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_226, A2 => lbl2_hscr_n_64, ZN => lbl2_hscr_n_251);
  lbl2_hscr_g18763 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_230, A2 => lbl2_hscr_n_3, ZN => lbl2_hscr_n_250);
  lbl2_hscr_g18764 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_123, A2 => lbl2_hscr_n_121, B => lbl2_hscr_n_226, ZN => lbl2_hscr_n_241);
  lbl2_hscr_g18765 : OA221D0BWP7T port map(A1 => lbl2_hscr_n_117, A2 => lbl2_hscr_n_12, B1 => lbl2_hscr_n_1, B2 => lbl2_hscr_n_141, C => lbl2_hscr_n_188, Z => lbl2_hscr_n_240);
  lbl2_hscr_g18766 : OAI31D0BWP7T port map(A1 => lbl2_hscr_n_64, A2 => lbl2_hscr_n_172, A3 => lbl2_hscr_n_174, B => lbl2_hscr_n_206, ZN => lbl2_hscr_n_239);
  lbl2_hscr_g18767 : OAI211D1BWP7T port map(A1 => lbl2_v_count(2), A2 => lbl2_hscr_n_30, B => lbl2_hscr_n_189, C => lbl2_hscr_n_151, ZN => lbl2_hscr_n_238);
  lbl2_hscr_g18768 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_55, A2 => lbl2_hscr_n_54, B => lbl2_hscr_n_205, C => lbl2_hscr_n_172, ZN => lbl2_hscr_n_246);
  lbl2_hscr_g18769 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_160, A2 => lbl2_hscr_n_133, A3 => lbl2_hscr_n_145, B1 => lbl2_hscr_n_202, B2 => lbl2_hscr_n_98, ZN => lbl2_hscr_n_245);
  lbl2_hscr_g18770 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_204, A2 => lbl2_hscr_n_172, A3 => lbl2_hscr_n_50, ZN => lbl2_hscr_n_244);
  lbl2_hscr_g18771 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_195, A2 => lbl2_v_count(1), A3 => lbl2_v_count(0), ZN => lbl2_hscr_n_243);
  lbl2_hscr_g18772 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_195, A2 => lbl2_hscr_n_116, A3 => lbl2_hscr_n_13, ZN => lbl2_hscr_n_242);
  lbl2_hscr_g18773 : CKND1BWP7T port map(I => lbl2_hscr_n_0, ZN => lbl2_hscr_n_237);
  lbl2_hscr_g18774 : INVD1BWP7T port map(I => lbl2_hscr_n_228, ZN => lbl2_hscr_n_227);
  lbl2_hscr_g18775 : OAI221D0BWP7T port map(A1 => lbl2_hscr_n_158, A2 => lbl2_hscr_n_64, B1 => lbl2_v_count(0), B2 => lbl2_hscr_n_99, C => lbl2_hscr_n_117, ZN => lbl2_hscr_n_225);
  lbl2_hscr_g18776 : NR2D0BWP7T port map(A1 => lbl2_hscr_n_193, A2 => lbl2_hscr_n_123, ZN => lbl2_hscr_n_224);
  lbl2_hscr_g18778 : AN2D0BWP7T port map(A1 => lbl2_hscr_n_205, A2 => lbl2_hscr_n_171, Z => lbl2_hscr_n_236);
  lbl2_hscr_g18779 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_117, B1 => lbl2_hscr_n_194, ZN => lbl2_hscr_n_235);
  lbl2_hscr_g18780 : NR2D0BWP7T port map(A1 => lbl2_hscr_n_193, A2 => lbl2_hscr_n_139, ZN => lbl2_hscr_n_234);
  lbl2_hscr_g18781 : OR2D1BWP7T port map(A1 => lbl2_hscr_n_197, A2 => lbl2_hscr_n_68, Z => lbl2_hscr_n_233);
  lbl2_hscr_g18782 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_193, A2 => lbl2_hscr_n_68, ZN => lbl2_hscr_n_232);
  lbl2_hscr_g18783 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_194, A2 => lbl2_v_count(0), ZN => lbl2_hscr_n_231);
  lbl2_hscr_g18784 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_194, A2 => lbl2_hscr_n_64, ZN => lbl2_hscr_n_230);
  lbl2_hscr_g18785 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_194, A2 => lbl2_v_count(1), ZN => lbl2_hscr_n_229);
  lbl2_hscr_g18786 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_194, A2 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_228);
  lbl2_hscr_g18787 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_196, A2 => lbl2_hscr_n_145, ZN => lbl2_hscr_n_226);
  lbl2_hscr_g18788 : OAI211D1BWP7T port map(A1 => lbl2_h_count(3), A2 => lbl2_hscr_n_45, B => lbl2_hscr_n_179, C => lbl2_hscr_n_88, ZN => lbl2_hscr_n_219);
  lbl2_hscr_g18789 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_80, A2 => lbl2_hscr_n_55, B => lbl2_hscr_n_194, ZN => lbl2_hscr_n_218);
  lbl2_hscr_g18790 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_76, A2 => lbl2_hscr_n_80, B => lbl2_hscr_n_204, ZN => lbl2_hscr_n_217);
  lbl2_hscr_g18791 : AO21D0BWP7T port map(A1 => lbl2_hscr_n_172, A2 => lbl2_hscr_n_80, B => lbl2_hscr_n_108, Z => lbl2_hscr_n_216);
  lbl2_hscr_g18792 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_133, A2 => lbl2_hscr_n_118, B => lbl2_hscr_n_202, ZN => lbl2_hscr_n_215);
  lbl2_hscr_g18793 : OR3XD1BWP7T port map(A1 => lbl2_hscr_n_104, A2 => lbl2_hscr_n_155, A3 => lbl2_hscr_n_193, Z => lbl2_hscr_n_214);
  lbl2_hscr_g18794 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_104, B1 => lbl2_hscr_n_172, B2 => lbl2_hscr_n_183, ZN => lbl2_hscr_n_213);
  lbl2_hscr_g18795 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_176, A2 => lbl2_hscr_n_162, B => lbl2_hscr_n_199, ZN => lbl2_hscr_n_212);
  lbl2_hscr_g18796 : AO21D0BWP7T port map(A1 => lbl2_hscr_n_158, A2 => lbl2_hscr_n_142, B => lbl2_hscr_n_207, Z => lbl2_hscr_n_211);
  lbl2_hscr_g18797 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_182, A2 => lbl2_hscr_n_120, A3 => lbl2_hscr_n_67, ZN => lbl2_hscr_n_223);
  lbl2_hscr_g18798 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_120, A2 => lbl2_hscr_n_98, B => lbl2_hscr_n_194, ZN => lbl2_hscr_n_222);
  lbl2_hscr_g18799 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_180, A2 => lbl2_hscr_n_132, A3 => lbl2_hscr_n_172, ZN => lbl2_hscr_n_221);
  lbl2_hscr_g18800 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_173, B1 => lbl2_hscr_n_82, B2 => lbl2_hscr_n_116, ZN => lbl2_hscr_n_220);
  lbl2_hscr_g18801 : INVD1BWP7T port map(I => lbl2_hscr_n_201, ZN => lbl2_hscr_n_202);
  lbl2_hscr_g18802 : INVD1BWP7T port map(I => lbl2_hscr_n_200, ZN => lbl2_hscr_n_199);
  lbl2_hscr_g18803 : INR2D1BWP7T port map(A1 => lbl2_hscr_n_183, B1 => lbl2_hscr_n_138, ZN => lbl2_hscr_n_210);
  lbl2_hscr_g18804 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_186, A2 => lbl2_h_count(2), ZN => lbl2_hscr_n_209);
  lbl2_hscr_g18805 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_182, A2 => lbl2_hscr_n_3, ZN => lbl2_hscr_n_208);
  lbl2_hscr_g18806 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_186, A2 => lbl2_hscr_n_3, ZN => lbl2_hscr_n_207);
  lbl2_hscr_g18807 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_175, A2 => lbl2_hscr_n_159, ZN => lbl2_hscr_n_206);
  lbl2_hscr_g18808 : INR2D1BWP7T port map(A1 => lbl2_hscr_n_180, B1 => lbl2_hscr_n_132, ZN => lbl2_hscr_n_205);
  lbl2_hscr_g18809 : AN2D1BWP7T port map(A1 => lbl2_hscr_n_180, A2 => lbl2_hscr_n_132, Z => lbl2_hscr_n_204);
  lbl2_hscr_g18810 : INR2XD0BWP7T port map(A1 => lbl2_hscr_n_92, B1 => lbl2_hscr_n_185, ZN => lbl2_hscr_n_203);
  lbl2_hscr_g18811 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_160, A2 => lbl2_hscr_n_172, ZN => lbl2_hscr_n_201);
  lbl2_hscr_g18812 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_183, A2 => lbl2_hscr_n_103, ZN => lbl2_hscr_n_200);
  lbl2_hscr_g18814 : INVD1BWP7T port map(I => lbl2_hscr_n_194, ZN => lbl2_hscr_n_193);
  lbl2_hscr_g18815 : AO31D1BWP7T port map(A1 => lbl2_hscr_n_145, A2 => lbl2_hscr_n_76, A3 => lbl2_hscr_n_48, B => lbl2_hscr_n_165, Z => lbl2_hscr_n_192);
  lbl2_hscr_g18816 : MOAI22D0BWP7T port map(A1 => lbl2_hscr_n_132, A2 => lbl2_hscr_n_134, B1 => lbl2_hscr_n_146, B2 => lbl2_hscr_n_160, ZN => lbl2_hscr_n_191);
  lbl2_hscr_g18817 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_161, B1 => lbl2_hscr_n_118, B2 => lbl2_hscr_n_160, ZN => lbl2_hscr_n_190);
  lbl2_hscr_g18818 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_39, A2 => lbl2_hscr_n_27, A3 => lbl2_v_count(2), B => lbl2_hscr_n_166, ZN => lbl2_hscr_n_189);
  lbl2_hscr_g18819 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_157, A2 => lbl2_hscr_n_98, B => lbl2_hscr_n_3, ZN => lbl2_hscr_n_188);
  lbl2_hscr_g18820 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_99, A2 => lbl2_hscr_n_46, B => lbl2_hscr_n_181, ZN => lbl2_hscr_n_187);
  lbl2_hscr_g18821 : NR2D0BWP7T port map(A1 => lbl2_hscr_n_171, A2 => lbl2_hscr_n_64, ZN => lbl2_hscr_n_198);
  lbl2_hscr_g18822 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_135, B1 => lbl2_hscr_n_172, B2 => lbl2_hscr_n_153, ZN => lbl2_hscr_n_197);
  lbl2_hscr_g18823 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_132, A2 => lbl2_hscr_n_171, ZN => lbl2_hscr_n_196);
  lbl2_hscr_g18824 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_131, A2 => lbl2_hscr_n_171, A3 => lbl2_hscr_n_104, ZN => lbl2_hscr_n_195);
  lbl2_hscr_g18825 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_131, A2 => lbl2_hscr_n_172, ZN => lbl2_hscr_n_194);
  lbl2_hscr_g18826 : INVD0BWP7T port map(I => lbl2_hscr_n_182, ZN => lbl2_hscr_n_181);
  lbl2_hscr_g18827 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_70, A2 => lbl2_hscr_n_19, A3 => lbl2_hscr_n_9, B => lbl2_hscr_n_400, ZN => lbl2_hscr_n_179);
  lbl2_hscr_g18828 : OR2D1BWP7T port map(A1 => lbl2_hscr_n_162, A2 => lbl2_hscr_n_120, Z => lbl2_hscr_n_178);
  lbl2_hscr_g18829 : IND3D1BWP7T port map(A1 => lbl2_central_x_vec(7), B1 => lbl2_hscr_n_29, B2 => lbl2_hscr_n_136, ZN => lbl2_hscr_n_177);
  lbl2_hscr_g18830 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_154, A2 => lbl2_hscr_n_101, ZN => lbl2_hscr_n_186);
  lbl2_hscr_g18831 : OAI211D1BWP7T port map(A1 => lbl2_n_124, A2 => lbl2_hscr_n_63, B => lbl2_hscr_n_136, C => lbl2_hscr_n_32, ZN => lbl2_hscr_n_185);
  lbl2_hscr_g18832 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_157, A2 => lbl2_hscr_n_131, ZN => lbl2_hscr_n_184);
  lbl2_hscr_g18833 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_154, A2 => lbl2_hscr_n_48, ZN => lbl2_hscr_n_183);
  lbl2_hscr_g18834 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_154, A2 => lbl2_hscr_n_82, ZN => lbl2_hscr_n_182);
  lbl2_hscr_g18835 : AOI211XD0BWP7T port map(A1 => lbl2_hscr_n_105, A2 => lbl2_central_x_vec(8), B => lbl2_hscr_n_129, C => lbl2_hscr_n_31, ZN => lbl2_hscr_n_180);
  lbl2_hscr_g18836 : INVD0BWP7T port map(I => lbl2_hscr_n_175, ZN => lbl2_hscr_n_174);
  lbl2_hscr_g18837 : INVD1BWP7T port map(I => lbl2_hscr_n_172, ZN => lbl2_hscr_n_171);
  lbl2_hscr_g18838 : MAOI22D0BWP7T port map(A1 => lbl2_hscr_n_47, A2 => lbl2_hscr_n_53, B1 => lbl2_hscr_n_143, B2 => lbl2_hscr_n_64, ZN => lbl2_hscr_n_170);
  lbl2_hscr_g18839 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_117, A2 => lbl2_v_count(1), B => lbl2_hscr_n_158, ZN => lbl2_hscr_n_169);
  lbl2_hscr_g18840 : AO21D0BWP7T port map(A1 => lbl2_hscr_n_133, A2 => lbl2_hscr_n_82, B => lbl2_hscr_n_163, Z => lbl2_hscr_n_168);
  lbl2_hscr_g18841 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_138, A2 => lbl2_hscr_n_2, B => lbl2_hscr_n_164, ZN => lbl2_hscr_n_167);
  lbl2_hscr_g18842 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_39, A2 => lbl2_hscr_n_130, B => lbl2_hscr_n_113, C => lbl2_hscr_n_112, ZN => lbl2_hscr_n_166);
  lbl2_hscr_g18843 : MOAI22D0BWP7T port map(A1 => lbl2_hscr_n_115, A2 => lbl2_hscr_n_145, B1 => lbl2_hscr_n_100, B2 => lbl2_hscr_n_50, ZN => lbl2_hscr_n_165);
  lbl2_hscr_g18844 : MOAI22D0BWP7T port map(A1 => lbl2_hscr_n_139, A2 => lbl2_hscr_n_2, B1 => lbl2_hscr_n_120, B2 => lbl2_hscr_n_13, ZN => lbl2_hscr_n_176);
  lbl2_hscr_g18845 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_131, A2 => lbl2_hscr_n_139, A3 => lbl2_v_count(0), ZN => lbl2_hscr_n_175);
  lbl2_hscr_g18846 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_133, A2 => lbl2_hscr_n_132, A3 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_173);
  lbl2_hscr_g18847 : MOAI22D1BWP7T port map(A1 => lbl2_hscr_n_109, A2 => lbl2_central_x_vec(6), B1 => lbl2_hscr_n_109, B2 => lbl2_central_x_vec(6), ZN => lbl2_hscr_n_172);
  lbl2_hscr_g18848 : INVD1BWP7T port map(I => lbl2_hscr_n_158, ZN => lbl2_hscr_n_157);
  lbl2_hscr_g18849 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_137, A2 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_164);
  lbl2_hscr_g18850 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_141, A2 => lbl2_v_count(1), ZN => lbl2_hscr_n_163);
  lbl2_hscr_g18851 : AN2D0BWP7T port map(A1 => lbl2_hscr_n_137, A2 => lbl2_v_count(0), Z => lbl2_hscr_n_162);
  lbl2_hscr_g18852 : NR2D0BWP7T port map(A1 => lbl2_hscr_n_101, A2 => lbl2_hscr_n_145, ZN => lbl2_hscr_n_156);
  lbl2_hscr_g18853 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_145, A2 => lbl2_hscr_n_82, ZN => lbl2_hscr_n_161);
  lbl2_hscr_g18854 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_132, A2 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_160);
  lbl2_hscr_g18855 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_145, A2 => lbl2_hscr_n_82, ZN => lbl2_hscr_n_159);
  lbl2_hscr_g18856 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_140, A2 => lbl2_v_count(0), ZN => lbl2_hscr_n_158);
  lbl2_hscr_g18857 : INVD0BWP7T port map(I => lbl2_hscr_n_154, ZN => lbl2_hscr_n_153);
  lbl2_hscr_g18859 : AOI33D1BWP7T port map(A1 => lbl2_hscr_n_72, A2 => lbl2_hscr_n_23, A3 => lbl2_hscr_n_1, B1 => lbl2_hscr_n_89, B2 => lbl2_h_count(1), B3 => lbl2_h_count(3), ZN => lbl2_hscr_n_151);
  lbl2_hscr_g18860 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_60, A2 => lbl2_hscr_n_70, B1 => lbl2_hscr_n_95, B2 => lbl2_v_count(1), C => lbl2_hscr_n_128, ZN => lbl2_hscr_n_150);
  lbl2_hscr_g18861 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_123, A2 => lbl2_v_count(0), B => lbl2_hscr_n_53, ZN => lbl2_hscr_n_149);
  lbl2_hscr_g18862 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_107, A2 => lbl2_hscr_n_13, B => lbl2_hscr_n_144, ZN => lbl2_hscr_n_148);
  lbl2_hscr_g18863 : OA21D0BWP7T port map(A1 => lbl2_hscr_n_125, A2 => lbl2_hscr_n_2, B => lbl2_hscr_n_134, Z => lbl2_hscr_n_147);
  lbl2_hscr_g18864 : OAI211D1BWP7T port map(A1 => lbl2_v_count(1), A2 => lbl2_hscr_n_99, B => lbl2_hscr_n_121, C => lbl2_hscr_n_96, ZN => lbl2_hscr_n_146);
  lbl2_hscr_g18865 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_90, B1 => lbl2_hscr_n_145, ZN => lbl2_hscr_n_155);
  lbl2_hscr_g18866 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_132, A2 => lbl2_hscr_n_116, ZN => lbl2_hscr_n_154);
  lbl2_hscr_g18867 : INVD1BWP7T port map(I => lbl2_hscr_n_116, ZN => lbl2_hscr_n_145);
  lbl2_hscr_g18868 : INR2D1BWP7T port map(A1 => lbl2_hscr_n_118, B1 => lbl2_hscr_n_13, ZN => lbl2_hscr_n_144);
  lbl2_hscr_g18869 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_120, A2 => lbl2_hscr_n_1, ZN => lbl2_hscr_n_143);
  lbl2_hscr_g18870 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_122, A2 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_142);
  lbl2_hscr_g18871 : OR2D1BWP7T port map(A1 => lbl2_hscr_n_117, A2 => lbl2_hscr_n_2, Z => lbl2_hscr_n_141);
  lbl2_hscr_g18872 : AN2D1BWP7T port map(A1 => lbl2_hscr_n_118, A2 => lbl2_hscr_n_1, Z => lbl2_hscr_n_140);
  lbl2_hscr_g18873 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_118, A2 => lbl2_v_count(1), ZN => lbl2_hscr_n_139);
  lbl2_hscr_g18874 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_122, A2 => lbl2_v_count(1), ZN => lbl2_hscr_n_138);
  lbl2_hscr_g18875 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_121, A2 => lbl2_v_count(1), ZN => lbl2_hscr_n_137);
  lbl2_hscr_g18876 : INVD1BWP7T port map(I => lbl2_hscr_n_134, ZN => lbl2_hscr_n_133);
  lbl2_hscr_g18877 : INVD1BWP7T port map(I => lbl2_hscr_n_132, ZN => lbl2_hscr_n_131);
  lbl2_hscr_g18878 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_86, A2 => lbl2_h_count(3), B1 => lbl2_hscr_n_27, B2 => FE_DBTN0_lbl2_v_count_2, ZN => lbl2_hscr_n_130);
  lbl2_hscr_g18879 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_105, A2 => lbl2_central_x_vec(8), A3 => lbl2_central_x_vec(7), ZN => lbl2_hscr_n_129);
  lbl2_hscr_g18880 : OAI33D1BWP7T port map(A1 => lbl2_v_count(0), A2 => lbl2_hscr_n_33, A3 => lbl2_hscr_n_81, B1 => lbl2_v_count(2), B2 => lbl2_hscr_n_36, B3 => lbl2_hscr_n_74, ZN => lbl2_hscr_n_128);
  lbl2_hscr_g18881 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_97, A2 => lbl2_v_count(1), B => lbl2_hscr_n_120, ZN => lbl2_hscr_n_127);
  lbl2_hscr_g18882 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_77, A2 => lbl2_hscr_n_17, A3 => lbl2_h_count(1), B1 => lbl2_hscr_n_85, B2 => lbl2_hscr_n_29, ZN => lbl2_hscr_n_126);
  lbl2_hscr_g18883 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_87, A2 => lbl2_hscr_n_78, A3 => lbl2_hscr_n_35, ZN => lbl2_hscr_n_136);
  lbl2_hscr_g18884 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_104, B1 => lbl2_hscr_n_1, B2 => lbl2_hscr_n_65, ZN => lbl2_hscr_n_135);
  lbl2_hscr_g18885 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_107, A2 => lbl2_hscr_n_83, A3 => lbl2_v_count(1), ZN => lbl2_hscr_n_134);
  lbl2_hscr_g18886 : MOAI22D1BWP7T port map(A1 => lbl2_hscr_n_105, A2 => lbl2_central_x_vec(7), B1 => lbl2_hscr_n_105, B2 => lbl2_central_x_vec(7), ZN => lbl2_hscr_n_132);
  lbl2_hscr_g18887 : INVD1BWP7T port map(I => lbl2_hscr_n_122, ZN => lbl2_hscr_n_121);
  lbl2_hscr_g18888 : INVD1BWP7T port map(I => lbl2_hscr_n_119, ZN => lbl2_hscr_n_120);
  lbl2_hscr_g18889 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_98, A2 => lbl2_hscr_n_97, ZN => lbl2_hscr_n_125);
  lbl2_hscr_g18890 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_97, A2 => lbl2_hscr_n_48, ZN => lbl2_hscr_n_124);
  lbl2_hscr_g18891 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_98, A2 => lbl2_v_count(1), ZN => lbl2_hscr_n_123);
  lbl2_hscr_g18892 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_99, A2 => lbl2_hscr_n_41, ZN => lbl2_hscr_n_122);
  lbl2_hscr_g18893 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_97, A2 => lbl2_hscr_n_41, ZN => lbl2_hscr_n_119);
  lbl2_hscr_g18894 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_96, A2 => lbl2_hscr_n_41, ZN => lbl2_hscr_n_118);
  lbl2_hscr_g18895 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_98, A2 => lbl2_hscr_n_41, ZN => lbl2_hscr_n_117);
  lbl2_hscr_g18896 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_50, A2 => lbl2_hscr_n_47, A3 => lbl2_v_count(3), B => lbl2_hscr_n_25, ZN => lbl2_hscr_n_115);
  lbl2_hscr_g18897 : AO21D0BWP7T port map(A1 => lbl2_hscr_n_82, A2 => lbl2_hscr_n_50, B => lbl2_hscr_n_54, Z => lbl2_hscr_n_114);
  lbl2_hscr_g18898 : OAI211D1BWP7T port map(A1 => FE_DBTN0_lbl2_v_count_2, A2 => lbl2_hscr_n_15, B => lbl2_hscr_n_77, C => lbl2_h_count(1), ZN => lbl2_hscr_n_113);
  lbl2_hscr_g18899 : IND4D0BWP7T port map(A1 => lbl2_hscr_n_62, B1 => lbl2_v_count(1), B2 => lbl2_hscr_n_14, B3 => lbl2_hscr_n_40, ZN => lbl2_hscr_n_112);
  lbl2_hscr_g18900 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_34, A2 => lbl2_hscr_n_13, A3 => lbl2_hscr_n_15, B1 => lbl2_hscr_n_401, B2 => lbl2_hscr_n_18, ZN => lbl2_hscr_n_111);
  lbl2_hscr_g18901 : OAI31D0BWP7T port map(A1 => lbl2_v_count(6), A2 => lbl2_v_count(2), A3 => lbl2_hscr_n_12, B => lbl2_hscr_n_93, ZN => lbl2_hscr_n_110);
  lbl2_hscr_g18902 : MAOI22D1BWP7T port map(A1 => lbl2_hscr_n_49, A2 => lbl2_central_x_vec(5), B1 => lbl2_hscr_n_49, B2 => lbl2_central_x_vec(5), ZN => lbl2_hscr_n_116);
  lbl2_hscr_g18903 : INVD0BWP7T port map(I => lbl2_hscr_n_107, ZN => lbl2_hscr_n_106);
  lbl2_hscr_g18904 : INVD0BWP7T port map(I => lbl2_hscr_n_103, ZN => lbl2_hscr_n_102);
  lbl2_hscr_g18905 : INVD0BWP7T port map(I => lbl2_hscr_n_101, ZN => lbl2_hscr_n_100);
  lbl2_hscr_g18906 : INVD1BWP7T port map(I => lbl2_hscr_n_99, ZN => lbl2_hscr_n_98);
  lbl2_hscr_g18907 : INVD1BWP7T port map(I => lbl2_hscr_n_97, ZN => lbl2_hscr_n_96);
  lbl2_hscr_g18908 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_49, B1 => lbl2_central_x_vec(5), ZN => lbl2_hscr_n_109);
  lbl2_hscr_g18909 : AN2D1BWP7T port map(A1 => lbl2_hscr_n_76, A2 => lbl2_v_count(3), Z => lbl2_hscr_n_108);
  lbl2_hscr_g18910 : INR2D1BWP7T port map(A1 => lbl2_hscr_n_41, B1 => lbl2_hscr_n_79, ZN => lbl2_hscr_n_107);
  lbl2_hscr_g18911 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_22, A2 => lbl2_hscr_n_49, ZN => lbl2_hscr_n_105);
  lbl2_hscr_g18912 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_41, B1 => lbl2_hscr_n_79, ZN => lbl2_hscr_n_104);
  lbl2_hscr_g18913 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_64, A2 => lbl2_h_count(2), ZN => lbl2_hscr_n_103);
  lbl2_hscr_g18914 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_64, A2 => lbl2_hscr_n_48, ZN => lbl2_hscr_n_101);
  lbl2_hscr_g18915 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_79, A2 => lbl2_hscr_n_83, ZN => lbl2_hscr_n_99);
  lbl2_hscr_g18916 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_79, A2 => lbl2_hscr_n_83, ZN => lbl2_hscr_n_97);
  lbl2_hscr_g18917 : INVD0BWP7T port map(I => lbl2_hscr_n_94, ZN => lbl2_hscr_n_95);
  lbl2_hscr_g18918 : CKND1BWP7T port map(I => lbl2_hscr_n_92, ZN => lbl2_hscr_n_93);
  lbl2_hscr_g18919 : MOAI22D0BWP7T port map(A1 => lbl2_hscr_n_14, A2 => lbl2_hscr_n_1, B1 => lbl2_hscr_n_39, B2 => lbl2_hscr_n_18, ZN => lbl2_hscr_n_89);
  lbl2_hscr_g18920 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_70, A2 => lbl2_hscr_n_42, B1 => lbl2_hscr_n_61, B2 => lbl2_hscr_n_29, ZN => lbl2_hscr_n_88);
  lbl2_hscr_g18921 : AOI211XD0BWP7T port map(A1 => lbl2_hscr_n_44, A2 => lbl2_h_count(3), B => lbl2_central_x_vec(8), C => lbl2_central_x_vec(7), ZN => lbl2_hscr_n_87);
  lbl2_hscr_g18922 : OAI31D0BWP7T port map(A1 => FE_DBTN1_lbl2_h_count_1, A2 => FE_DBTN0_lbl2_v_count_2, A3 => lbl2_hscr_n_43, B => lbl2_hscr_n_14, ZN => lbl2_hscr_n_86);
  lbl2_hscr_g18923 : IOA21D0BWP7T port map(A1 => lbl2_hscr_n_18, A2 => lbl2_v_count(0), B => lbl2_hscr_n_45, ZN => lbl2_hscr_n_85);
  lbl2_hscr_g18924 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_11, A2 => lbl2_hscr_n_37, A3 => lbl2_h_count(1), B1 => lbl2_hscr_n_70, B2 => lbl2_hscr_n_13, ZN => lbl2_hscr_n_84);
  lbl2_hscr_g18925 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_21, B1 => lbl2_v_count(0), B2 => lbl2_hscr_n_72, ZN => lbl2_hscr_n_94);
  lbl2_hscr_g18926 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_73, A2 => lbl2_v_count(7), A3 => lbl2_v_count(8), ZN => lbl2_hscr_n_92);
  lbl2_hscr_g18927 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_64, A2 => lbl2_hscr_n_47, ZN => lbl2_hscr_n_91);
  lbl2_hscr_g18928 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_82, A2 => lbl2_hscr_n_48, ZN => lbl2_hscr_n_90);
  lbl2_hscr_g18929 : INVD1BWP7T port map(I => lbl2_hscr_n_65, ZN => lbl2_hscr_n_83);
  lbl2_hscr_g18930 : INVD1BWP7T port map(I => lbl2_hscr_n_64, ZN => lbl2_hscr_n_82);
  lbl2_hscr_g18931 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_54, A2 => lbl2_hscr_n_10, B => lbl2_v_count(8), ZN => lbl2_hscr_n_78);
  lbl2_hscr_g18932 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_42, B1 => lbl2_hscr_n_72, ZN => lbl2_hscr_n_81);
  lbl2_hscr_g18933 : INR2D1BWP7T port map(A1 => lbl2_hscr_n_50, B1 => lbl2_v_count(3), ZN => lbl2_hscr_n_80);
  lbl2_hscr_g18934 : OA211D0BWP7T port map(A1 => lbl2_v_count(4), A2 => lbl2_hscr_n_17, B => lbl2_hscr_n_46, C => lbl2_hscr_n_30, Z => lbl2_hscr_n_79);
  lbl2_hscr_g18936 : OA21D0BWP7T port map(A1 => lbl2_hscr_n_43, A2 => FE_DBTN1_lbl2_h_count_1, B => lbl2_hscr_n_40, Z => lbl2_hscr_n_74);
  lbl2_hscr_g18937 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_40, A2 => lbl2_hscr_n_21, A3 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_77);
  lbl2_hscr_g18938 : AN3D1BWP7T port map(A1 => lbl2_hscr_n_50, A2 => lbl2_hscr_n_30, A3 => lbl2_hscr_n_26, Z => lbl2_hscr_n_76);
  lbl2_hscr_g18939 : INVD0BWP7T port map(I => lbl2_hscr_n_68, ZN => lbl2_hscr_n_67);
  lbl2_hscr_g18940 : AOI211D1BWP7T port map(A1 => lbl2_central_x_vec(5), A2 => lbl2_h_count(4), B => lbl2_hscr_n_20, C => lbl2_hscr_n_24, ZN => lbl2_hscr_n_66);
  lbl2_hscr_g18941 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_52, A2 => lbl2_hscr_n_10, ZN => lbl2_hscr_n_73);
  lbl2_hscr_g18942 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_56, A2 => lbl2_hscr_n_40, ZN => lbl2_hscr_n_72);
  lbl2_hscr_g18943 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_48, A2 => lbl2_h_count(2), ZN => lbl2_hscr_n_71);
  lbl2_hscr_g18944 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_57, A2 => lbl2_hscr_n_39, ZN => lbl2_hscr_n_70);
  lbl2_hscr_g18946 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_47, A2 => lbl2_h_count(2), ZN => lbl2_hscr_n_68);
  lbl2_hscr_g18947 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_22, A2 => FE_DBTN2_lbl2_h_count_3, B => lbl2_hscr_n_44, ZN => lbl2_hscr_n_63);
  lbl2_hscr_g18948 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_34, A2 => lbl2_v_count(0), B => lbl2_hscr_n_23, ZN => lbl2_hscr_n_62);
  lbl2_hscr_g18949 : MOAI22D0BWP7T port map(A1 => lbl2_hscr_n_12, A2 => lbl2_h_count(3), B1 => lbl2_hscr_n_19, B2 => lbl2_v_count(1), ZN => lbl2_hscr_n_61);
  lbl2_hscr_g18950 : MOAI22D0BWP7T port map(A1 => lbl2_hscr_n_12, A2 => lbl2_hscr_n_21, B1 => lbl2_hscr_n_29, B2 => lbl2_hscr_n_19, ZN => lbl2_hscr_n_60);
  lbl2_hscr_g18951 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_35, A2 => lbl2_v_count(5), B => lbl2_v_count(4), ZN => lbl2_hscr_n_59);
  lbl2_hscr_g18952 : MOAI22D0BWP7T port map(A1 => lbl2_central_x_vec(7), A2 => lbl2_hscr_n_20, B1 => lbl2_central_x_vec(6), B2 => lbl2_hscr_n_20, ZN => lbl2_hscr_n_58);
  lbl2_hscr_g18953 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_16, A2 => lbl2_v_count(3), B => lbl2_hscr_n_53, ZN => lbl2_hscr_n_65);
  lbl2_hscr_g18954 : AOI21D1BWP7T port map(A1 => lbl2_hscr_n_28, A2 => lbl2_h_count(4), B => lbl2_hscr_n_49, ZN => lbl2_hscr_n_64);
  lbl2_hscr_g18955 : INVD0BWP7T port map(I => lbl2_hscr_n_56, ZN => lbl2_hscr_n_57);
  lbl2_hscr_g18956 : INVD1BWP7T port map(I => lbl2_hscr_n_52, ZN => lbl2_hscr_n_51);
  lbl2_hscr_g18957 : INVD1BWP7T port map(I => lbl2_hscr_n_48, ZN => lbl2_hscr_n_47);
  lbl2_hscr_g18958 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_37, A2 => lbl2_hscr_n_15, ZN => lbl2_hscr_n_56);
  lbl2_hscr_g18959 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_26, A2 => lbl2_v_count(5), ZN => lbl2_hscr_n_55);
  lbl2_hscr_g18960 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_30, A2 => lbl2_v_count(5), ZN => lbl2_hscr_n_54);
  lbl2_hscr_g18961 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_16, A2 => lbl2_v_count(3), ZN => lbl2_hscr_n_53);
  lbl2_hscr_g18962 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_25, A2 => lbl2_v_count(5), ZN => lbl2_hscr_n_52);
  lbl2_hscr_g18963 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_26, A2 => lbl2_v_count(5), ZN => lbl2_hscr_n_50);
  lbl2_hscr_g18964 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_28, A2 => lbl2_h_count(4), ZN => lbl2_hscr_n_49);
  lbl2_hscr_g18965 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_28, A2 => lbl2_hscr_n_36, ZN => lbl2_hscr_n_48);
  lbl2_hscr_g18966 : INVD1BWP7T port map(I => lbl2_hscr_n_40, ZN => lbl2_hscr_n_39);
  lbl2_hscr_g18968 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_17, A2 => lbl2_hscr_n_25, ZN => lbl2_hscr_n_46);
  lbl2_hscr_g18969 : CKND2D0BWP7T port map(A1 => lbl2_hscr_n_11, A2 => lbl2_v_count(2), ZN => lbl2_hscr_n_45);
  lbl2_hscr_g18970 : INR2D1BWP7T port map(A1 => lbl2_h_count(4), B1 => lbl2_hscr_n_22, ZN => lbl2_hscr_n_44);
  lbl2_hscr_g18971 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_2, A2 => lbl2_h_count(0), B => lbl2_hscr_n_1, ZN => lbl2_hscr_n_43);
  lbl2_hscr_g18972 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_1, A2 => lbl2_h_count(1), B1 => lbl2_v_count(1), B2 => FE_DBTN1_lbl2_h_count_1, ZN => lbl2_hscr_n_42);
  lbl2_hscr_g18973 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_1, A2 => lbl2_v_count(2), B => lbl2_hscr_n_18, ZN => lbl2_hscr_n_41);
  lbl2_hscr_g18974 : MAOI22D0BWP7T port map(A1 => lbl2_v_count(2), A2 => lbl2_v_count(3), B1 => lbl2_v_count(2), B2 => lbl2_v_count(3), ZN => lbl2_hscr_n_40);
  lbl2_hscr_g18975 : INVD0BWP7T port map(I => lbl2_hscr_n_34, ZN => lbl2_hscr_n_33);
  lbl2_hscr_g18976 : INVD0BWP7T port map(I => lbl2_hscr_n_32, ZN => lbl2_hscr_n_31);
  lbl2_hscr_g18977 : INVD0BWP7T port map(I => lbl2_hscr_n_28, ZN => lbl2_hscr_n_27);
  lbl2_hscr_g18978 : INVD1BWP7T port map(I => lbl2_hscr_n_26, ZN => lbl2_hscr_n_25);
  lbl2_hscr_g18979 : NR2XD0BWP7T port map(A1 => lbl2_h_count(4), A2 => direction_in(2), ZN => lbl2_hscr_n_24);
  lbl2_hscr_g18980 : NR2D0BWP7T port map(A1 => lbl2_h_count(2), A2 => lbl2_v_count(2), ZN => lbl2_hscr_n_37);
  lbl2_hscr_g18981 : ND2D1BWP7T port map(A1 => lbl2_h_count(2), A2 => lbl2_h_count(3), ZN => lbl2_hscr_n_36);
  lbl2_hscr_g18982 : NR2XD0BWP7T port map(A1 => lbl2_v_count(7), A2 => lbl2_v_count(8), ZN => lbl2_hscr_n_35);
  lbl2_hscr_g18983 : NR2D0BWP7T port map(A1 => lbl2_h_count(3), A2 => lbl2_h_count(0), ZN => lbl2_hscr_n_34);
  lbl2_hscr_g18984 : ND2D1BWP7T port map(A1 => lbl2_central_x_vec(8), A2 => lbl2_central_x_vec(7), ZN => lbl2_hscr_n_32);
  lbl2_hscr_g18985 : OR2D1BWP7T port map(A1 => lbl2_v_count(3), A2 => lbl2_v_count(4), Z => lbl2_hscr_n_30);
  lbl2_hscr_g18986 : NR2D1BWP7T port map(A1 => lbl2_h_count(1), A2 => lbl2_h_count(0), ZN => lbl2_hscr_n_29);
  lbl2_hscr_g18987 : CKND2D1BWP7T port map(A1 => FE_DBTN2_lbl2_h_count_3, A2 => lbl2_hscr_n_3, ZN => lbl2_hscr_n_28);
  lbl2_hscr_g18988 : CKND2D1BWP7T port map(A1 => lbl2_v_count(4), A2 => lbl2_v_count(3), ZN => lbl2_hscr_n_26);
  lbl2_hscr_g18989 : INVD0BWP7T port map(I => lbl2_hscr_n_17, ZN => lbl2_hscr_n_16);
  lbl2_hscr_g18990 : INVD0BWP7T port map(I => lbl2_hscr_n_15, ZN => lbl2_hscr_n_14);
  lbl2_hscr_g18991 : INVD0BWP7T port map(I => lbl2_hscr_n_12, ZN => lbl2_hscr_n_11);
  lbl2_hscr_g18992 : NR2D0BWP7T port map(A1 => lbl2_h_count(3), A2 => lbl2_h_count(1), ZN => lbl2_hscr_n_23);
  lbl2_hscr_g18993 : ND2D1BWP7T port map(A1 => lbl2_central_x_vec(6), A2 => lbl2_central_x_vec(5), ZN => lbl2_hscr_n_22);
  lbl2_hscr_g18994 : ND2D1BWP7T port map(A1 => lbl2_h_count(3), A2 => lbl2_h_count(0), ZN => lbl2_hscr_n_21);
  lbl2_hscr_g18995 : NR2XD0BWP7T port map(A1 => lbl2_central_x_vec(5), A2 => lbl2_h_count(4), ZN => lbl2_hscr_n_20);
  lbl2_hscr_g18996 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_2, A2 => lbl2_h_count(3), ZN => lbl2_hscr_n_19);
  lbl2_hscr_g18997 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_1, A2 => lbl2_v_count(2), ZN => lbl2_hscr_n_18);
  lbl2_hscr_g18998 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_1, A2 => FE_DBTN0_lbl2_v_count_2, ZN => lbl2_hscr_n_17);
  lbl2_hscr_g18999 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_3, A2 => FE_DBTN0_lbl2_v_count_2, ZN => lbl2_hscr_n_15);
  lbl2_hscr_g19000 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_1, A2 => lbl2_v_count(0), ZN => lbl2_hscr_n_13);
  lbl2_hscr_g19001 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_1, A2 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_12);
  lbl2_hscr_g19002 : INVD1BWP7T port map(I => lbl2_v_count(6), ZN => lbl2_hscr_n_10);
  lbl2_hscr_g19003 : INVD1BWP7T port map(I => lbl2_h_count(0), ZN => lbl2_hscr_n_9);
  lbl2_hscr_g19006 : INVD0BWP7T port map(I => lbl2_central_x_vec(6), ZN => lbl2_hscr_n_6);
  lbl2_hscr_g19009 : INVD1BWP7T port map(I => lbl2_h_count(2), ZN => lbl2_hscr_n_3);
  lbl2_hscr_g19010 : INVD1BWP7T port map(I => lbl2_v_count(0), ZN => lbl2_hscr_n_2);
  lbl2_hscr_g19011 : INVD1BWP7T port map(I => lbl2_v_count(1), ZN => lbl2_hscr_n_1);
  lbl2_hscr_g2 : INR2D1BWP7T port map(A1 => lbl2_hscr_n_196, B1 => lbl2_hscr_n_139, ZN => lbl2_hscr_n_0);
  lbl2_hscr_g19012 : INVD0BWP7T port map(I => lbl2_v_count(8), ZN => lbl2_hscr_n_38);
  lbl2_hscr_g19014 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_111, A2 => lbl2_hscr_n_40, B => lbl2_hscr_n_94, ZN => lbl2_hscr_n_400);
  lbl2_hscr_g19015 : AO21D0BWP7T port map(A1 => lbl2_hscr_n_27, A2 => lbl2_hscr_n_9, B => lbl2_hscr_n_19, Z => lbl2_hscr_n_401);
  lbl2_pxl_g8179 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_208, A2 => lbl2_pxl_n_191, A3 => lbl2_pxl_n_125, A4 => lbl2_pxl_n_104, ZN => lbl2_pixelator_color(2));
  lbl2_pxl_g8180 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_210, A2 => lbl2_pxl_n_191, A3 => lbl2_pxl_n_177, ZN => lbl2_pixelator_color(0));
  lbl2_pxl_g8181 : ND4D0BWP7T port map(A1 => lbl2_pxl_n_207, A2 => lbl2_pxl_n_184, A3 => lbl2_pxl_n_181, A4 => lbl2_pxl_n_185, ZN => lbl2_pxl_n_210);
  lbl2_pxl_g8182 : AN3D0BWP7T port map(A1 => lbl2_pxl_n_206, A2 => lbl2_pxl_n_195, A3 => lbl2_pxl_n_120, Z => lbl2_pixelator_color(3));
  lbl2_pxl_g8183 : ND4D0BWP7T port map(A1 => lbl2_pxl_n_205, A2 => lbl2_pxl_n_195, A3 => lbl2_pxl_n_167, A4 => lbl2_pxl_n_159, ZN => lbl2_pxl_n_208);
  lbl2_pxl_g8184 : AN4D0BWP7T port map(A1 => lbl2_pxl_n_201, A2 => lbl2_pxl_n_194, A3 => lbl2_pxl_n_197, A4 => lbl2_pxl_n_167, Z => lbl2_pxl_n_207);
  lbl2_pxl_g8185 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_203, A2 => lbl2_pxl_n_175, A3 => lbl2_pxl_n_125, ZN => lbl2_pxl_n_206);
  lbl2_pxl_g8186 : AOI211XD0BWP7T port map(A1 => lbl2_pxl_n_176, A2 => position_0(10), B => lbl2_pxl_n_202, C => lbl2_pxl_n_157, ZN => lbl2_pxl_n_205);
  lbl2_pxl_g8187 : AN4D1BWP7T port map(A1 => lbl2_pxl_n_199, A2 => lbl2_pxl_n_195, A3 => lbl2_pxl_n_198, A4 => lbl2_pxl_n_178, Z => lbl2_pixelator_color(1));
  lbl2_pxl_g8188 : ND4D0BWP7T port map(A1 => lbl2_pxl_n_199, A2 => lbl2_pxl_n_184, A3 => lbl2_pxl_n_179, A4 => lbl2_pxl_n_173, ZN => lbl2_pxl_n_203);
  lbl2_pxl_g8189 : OAI31D0BWP7T port map(A1 => lbl2_pxl_n_124, A2 => lbl2_pxl_n_136, A3 => lbl2_pxl_n_183, B => lbl2_pxl_n_200, ZN => lbl2_pxl_n_202);
  lbl2_pxl_g8190 : OA221D0BWP7T port map(A1 => lbl2_pxl_n_193, A2 => lbl2_pxl_n_163, B1 => lbl2_pxl_n_160, B2 => lbl2_pxl_n_187, C => lbl2_pxl_n_186, Z => lbl2_pxl_n_201);
  lbl2_pxl_g8191 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_196, A2 => lbl2_pxl_n_188, A3 => lbl2_pxl_n_180, A4 => lbl2_pxl_n_177, ZN => lbl2_pxl_n_200);
  lbl2_pxl_g8192 : IINR4D0BWP7T port map(A1 => lbl2_pxl_n_181, A2 => lbl2_pxl_n_2, B1 => lbl2_pxl_n_190, B2 => lbl2_pxl_n_180, ZN => lbl2_pxl_n_198);
  lbl2_pxl_g8193 : OA21D0BWP7T port map(A1 => lbl2_pxl_n_193, A2 => lbl2_pxl_n_155, B => lbl2_pxl_n_194, Z => lbl2_pxl_n_199);
  lbl2_pxl_g8194 : IINR4D0BWP7T port map(A1 => lbl2_pxl_n_158, A2 => lbl2_pxl_n_120, B1 => lbl2_pxl_n_189, B2 => lbl2_pxl_n_104, ZN => lbl2_pxl_n_197);
  lbl2_pxl_g8195 : OAI22D0BWP7T port map(A1 => lbl2_pxl_n_193, A2 => lbl2_pxl_n_164, B1 => lbl2_pxl_n_187, B2 => lbl2_pxl_n_149, ZN => lbl2_pxl_n_196);
  lbl2_pxl_g8196 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_193, B1 => lbl2_pxl_n_113, B2 => lbl2_pxl_n_148, ZN => lbl2_pxl_n_195);
  lbl2_pxl_g8197 : IND4D0BWP7T port map(A1 => lbl2_pxl_n_113, B1 => lbl2_pxl_n_116, B2 => lbl2_pxl_n_148, B3 => lbl2_pxl_n_192, ZN => lbl2_pxl_n_194);
  lbl2_pxl_g8198 : INVD1BWP7T port map(I => lbl2_pxl_n_192, ZN => lbl2_pxl_n_193);
  lbl2_pxl_g8199 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_187, A2 => lbl2_pxl_n_150, A3 => lbl2_pxl_n_131, ZN => lbl2_pxl_n_192);
  lbl2_pxl_g8200 : OAI211D1BWP7T port map(A1 => lbl2_pxl_n_88, A2 => lbl2_pxl_n_174, B => lbl2_pxl_n_158, C => lbl2_pxl_n_159, ZN => lbl2_pxl_n_190);
  lbl2_pxl_g8201 : IND4D0BWP7T port map(A1 => lbl2_pxl_n_175, B1 => lbl2_pxl_n_173, B2 => lbl2_pxl_n_178, B3 => lbl2_pxl_n_2, ZN => lbl2_pxl_n_191);
  lbl2_pxl_g8202 : OAI32D1BWP7T port map(A1 => lbl2_pxl_n_126, A2 => lbl2_pxl_n_123, A3 => lbl2_pxl_n_152, B1 => lbl2_pxl_n_111, B2 => lbl2_pxl_n_183, ZN => lbl2_pxl_n_189);
  lbl2_pxl_g8203 : OAI22D0BWP7T port map(A1 => lbl2_pxl_n_183, A2 => lbl2_pxl_n_107, B1 => lbl2_pxl_n_174, B2 => lbl2_pxl_n_112, ZN => lbl2_pxl_n_188);
  lbl2_pxl_g8204 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_183, B1 => lbl2_pxl_n_151, ZN => lbl2_pxl_n_187);
  lbl2_pxl_g8205 : IND4D0BWP7T port map(A1 => lbl2_pxl_n_124, B1 => lbl2_pxl_n_139, B2 => lbl2_pxl_n_136, B3 => lbl2_pxl_n_182, ZN => lbl2_pxl_n_186);
  lbl2_pxl_g8206 : AOI222D0BWP7T port map(A1 => lbl2_pxl_n_170, A2 => position_1(10), B1 => lbl2_pxl_n_165, B2 => lbl2_pxl_n_143, C1 => lbl2_pxl_n_169, C2 => lbl2_pxl_n_147, ZN => lbl2_pxl_n_185);
  lbl2_pxl_g8207 : INVD1BWP7T port map(I => lbl2_pxl_n_182, ZN => lbl2_pxl_n_183);
  lbl2_pxl_g8208 : OR2D1BWP7T port map(A1 => lbl2_pxl_n_174, A2 => lbl2_pxl_n_118, Z => lbl2_pxl_n_184);
  lbl2_pxl_g8209 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_174, A2 => lbl2_pxl_n_142, ZN => lbl2_pxl_n_182);
  lbl2_pxl_g8210 : AO21D0BWP7T port map(A1 => lbl2_pxl_n_112, A2 => lbl2_pxl_n_88, B => lbl2_pxl_n_174, Z => lbl2_pxl_n_179);
  lbl2_pxl_g8211 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_174, B1 => player_state_1(0), B2 => lbl2_pxl_n_115, ZN => lbl2_pxl_n_181);
  lbl2_pxl_g8212 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_174, A2 => lbl2_pxl_n_114, A3 => player_state_1(0), ZN => lbl2_pxl_n_180);
  lbl2_pxl_g8213 : OAI221D0BWP7T port map(A1 => lbl2_pxl_n_166, A2 => lbl2_pxl_n_127, B1 => lbl2_pxl_n_130, B2 => lbl2_pxl_n_161, C => lbl2_pxl_n_168, ZN => lbl2_pxl_n_176);
  lbl2_pxl_g8214 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_172, A2 => lbl2_pxl_n_119, ZN => lbl2_pxl_n_178);
  lbl2_pxl_g8215 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_171, A2 => lbl2_pxl_n_99, ZN => lbl2_pxl_n_177);
  lbl2_pxl_g8216 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_171, A2 => lbl2_pxl_n_119, A3 => lbl2_pxl_n_97, A4 => lbl2_data_synced(7), ZN => lbl2_pxl_n_175);
  lbl2_pxl_g8218 : IND4D0BWP7T port map(A1 => lbl2_pxl_n_119, B1 => lbl2_pxl_n_97, B2 => lbl2_pxl_n_99, B3 => lbl2_pxl_n_172, ZN => lbl2_pxl_n_174);
  lbl2_pxl_g8219 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_147, B1 => lbl2_pxl_n_121, B2 => lbl2_pxl_n_169, ZN => lbl2_pxl_n_173);
  lbl2_pxl_g8220 : INVD0BWP7T port map(I => lbl2_pxl_n_172, ZN => lbl2_pxl_n_171);
  lbl2_pxl_g8221 : OAI22D0BWP7T port map(A1 => lbl2_pxl_n_166, A2 => lbl2_pxl_n_132, B1 => lbl2_pxl_n_161, B2 => lbl2_pxl_n_138, ZN => lbl2_pxl_n_170);
  lbl2_pxl_g8222 : INR3D0BWP7T port map(A1 => lbl2_pxl_n_169, B1 => lbl2_pxl_n_121, B2 => lbl2_pxl_n_147, ZN => lbl2_pxl_n_172);
  lbl2_pxl_g8223 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_131, A2 => position_1(10), B1 => lbl2_pxl_n_128, B2 => position_0(10), C => lbl2_pxl_n_166, ZN => lbl2_pxl_n_169);
  lbl2_pxl_g8224 : AOI32D1BWP7T port map(A1 => lbl2_pxl_n_165, A2 => lbl2_pxl_n_144, A3 => lbl2_pxl_n_134, B1 => lbl2_pxl_n_156, B2 => lbl2_pxl_n_137, ZN => lbl2_pxl_n_168);
  lbl2_pxl_g8225 : IND4D0BWP7T port map(A1 => lbl2_pxl_n_155, B1 => lbl2_pxl_n_100, B2 => lbl2_pxl_n_132, B3 => lbl2_pxl_n_162, ZN => lbl2_pxl_n_167);
  lbl2_pxl_g8226 : OAI211D1BWP7T port map(A1 => lbl2_pxl_n_8, A2 => lbl2_pxl_n_135, B => lbl2_pxl_n_165, C => lbl2_pxl_n_144, ZN => lbl2_pxl_n_166);
  lbl2_pxl_g8227 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_129, A2 => position_0(10), B1 => lbl2_pxl_n_139, B2 => position_1(10), C => lbl2_pxl_n_161, ZN => lbl2_pxl_n_165);
  lbl2_pxl_g8228 : OA31D1BWP7T port map(A1 => lbl2_data_synced(3), A2 => lbl2_pxl_n_100, A3 => lbl2_pxl_n_155, B => lbl2_pxl_n_127, Z => lbl2_pxl_n_164);
  lbl2_pxl_g8229 : MAOI22D0BWP7T port map(A1 => lbl2_pxl_n_127, A2 => lbl2_pxl_n_140, B1 => lbl2_pxl_n_155, B2 => lbl2_pxl_n_106, ZN => lbl2_pxl_n_163);
  lbl2_pxl_g8230 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_154, A2 => lbl2_pxl_n_150, ZN => lbl2_pxl_n_162);
  lbl2_pxl_g8231 : MAOI22D0BWP7T port map(A1 => lbl2_pxl_n_130, A2 => lbl2_pxl_n_133, B1 => lbl2_pxl_n_150, B2 => lbl2_pxl_n_132, ZN => lbl2_pxl_n_160);
  lbl2_pxl_g8232 : OAI211D1BWP7T port map(A1 => lbl2_pxl_n_8, A2 => lbl2_pxl_n_136, B => lbl2_pxl_n_156, C => lbl2_pxl_n_141, ZN => lbl2_pxl_n_161);
  lbl2_pxl_g8233 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_152, A2 => lbl2_pxl_n_141, ZN => lbl2_pxl_n_157);
  lbl2_pxl_g8234 : IND2D1BWP7T port map(A1 => player_state_1(0), B1 => lbl2_pxl_n_153, ZN => lbl2_pxl_n_159);
  lbl2_pxl_g8235 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_153, A2 => player_state_1(0), ZN => lbl2_pxl_n_158);
  lbl2_pxl_g8236 : ND4D0BWP7T port map(A1 => lbl2_pxl_n_151, A2 => lbl2_pxl_n_122, A3 => lbl2_pxl_n_95, A4 => lbl2_pxl_n_87, ZN => lbl2_pxl_n_154);
  lbl2_pxl_g8237 : INR2XD0BWP7T port map(A1 => lbl2_pxl_n_123, B1 => lbl2_pxl_n_152, ZN => lbl2_pxl_n_156);
  lbl2_pxl_g8238 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_113, B1 => lbl2_pxl_n_117, B2 => lbl2_pxl_n_148, ZN => lbl2_pxl_n_155);
  lbl2_pxl_g8239 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_145, A2 => lbl2_pxl_n_109, ZN => lbl2_pxl_n_153);
  lbl2_pxl_g8240 : OAI211D1BWP7T port map(A1 => lbl2_pxl_n_94, A2 => lbl2_pxl_n_54, B => lbl2_pxl_n_146, C => lbl2_pxl_n_109, ZN => lbl2_pxl_n_152);
  lbl2_pxl_g8241 : OA21D0BWP7T port map(A1 => lbl2_pxl_n_135, A2 => lbl2_pxl_n_133, B => lbl2_pxl_n_130, Z => lbl2_pxl_n_149);
  lbl2_pxl_g8242 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_139, A2 => lbl2_pxl_n_137, A3 => lbl2_pxl_n_124, ZN => lbl2_pxl_n_151);
  lbl2_pxl_g8243 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_133, B1 => lbl2_pxl_n_135, B2 => lbl2_pxl_n_130, ZN => lbl2_pxl_n_150);
  lbl2_pxl_g8244 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_140, A2 => lbl2_pxl_n_128, ZN => lbl2_pxl_n_148);
  lbl2_pxl_g8245 : AN2D1BWP7T port map(A1 => lbl2_pxl_n_140, A2 => position_1(10), Z => lbl2_pxl_n_147);
  lbl2_pxl_g8246 : CKND1BWP7T port map(I => lbl2_pxl_n_145, ZN => lbl2_pxl_n_146);
  lbl2_pxl_g8247 : INVD0BWP7T port map(I => lbl2_pxl_n_144, ZN => lbl2_pxl_n_143);
  lbl2_pxl_g8248 : OAI211D1BWP7T port map(A1 => lbl2_pxl_n_111, A2 => lbl2_pxl_n_107, B => lbl2_pxl_n_122, C => lbl2_pxl_n_105, ZN => lbl2_pxl_n_142);
  lbl2_pxl_g8249 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_125, B1 => lbl2_pxl_n_91, B2 => lbl2_pxl_n_120, ZN => lbl2_pxl_n_145);
  lbl2_pxl_g8250 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_133, A2 => position_1(10), ZN => lbl2_pxl_n_144);
  lbl2_pxl_g8251 : INVD0BWP7T port map(I => lbl2_pxl_n_139, ZN => lbl2_pxl_n_138);
  lbl2_pxl_g8252 : INVD0BWP7T port map(I => lbl2_pxl_n_137, ZN => lbl2_pxl_n_136);
  lbl2_pxl_g8253 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_123, A2 => lbl2_pxl_n_126, ZN => lbl2_pxl_n_141);
  lbl2_pxl_g8254 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_108, A2 => lbl2_pxl_n_1, A3 => lbl2_pxl_n_30, ZN => lbl2_pxl_n_140);
  lbl2_pxl_g8255 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_1, A2 => lbl2_pxl_n_103, A3 => lbl2_pxl_n_6, A4 => lbl2_pxl_n_16, ZN => lbl2_pxl_n_139);
  lbl2_pxl_g8256 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_0, A2 => lbl2_pxl_n_103, A3 => lbl2_pxl_n_6, A4 => lbl2_pxl_n_23, ZN => lbl2_pxl_n_137);
  lbl2_pxl_g8257 : INVD0BWP7T port map(I => lbl2_pxl_n_135, ZN => lbl2_pxl_n_134);
  lbl2_pxl_g8258 : INVD1BWP7T port map(I => lbl2_pxl_n_132, ZN => lbl2_pxl_n_131);
  lbl2_pxl_g8259 : INVD1BWP7T port map(I => lbl2_pxl_n_129, ZN => lbl2_pxl_n_130);
  lbl2_pxl_g8260 : INVD0BWP7T port map(I => lbl2_pxl_n_128, ZN => lbl2_pxl_n_127);
  lbl2_pxl_g8261 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_0, B1 => lbl2_pxl_n_20, B2 => lbl2_pxl_n_110, ZN => lbl2_pxl_n_135);
  lbl2_pxl_g8262 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_1, A2 => lbl2_pxl_n_102, A3 => lbl2_dx(3), A4 => lbl2_pxl_n_29, ZN => lbl2_pxl_n_133);
  lbl2_pxl_g8263 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_1, B1 => lbl2_pxl_n_25, B2 => lbl2_pxl_n_110, ZN => lbl2_pxl_n_132);
  lbl2_pxl_g8264 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_0, A2 => lbl2_pxl_n_102, A3 => lbl2_dx(3), A4 => lbl2_pxl_n_27, ZN => lbl2_pxl_n_129);
  lbl2_pxl_g8265 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_108, A2 => lbl2_pxl_n_0, A3 => lbl2_pxl_n_18, ZN => lbl2_pxl_n_128);
  lbl2_pxl_g8266 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_107, A2 => lbl2_pxl_n_8, ZN => lbl2_pxl_n_126);
  lbl2_pxl_g8267 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_112, A2 => lbl2_pxl_n_8, ZN => lbl2_pxl_n_125);
  lbl2_pxl_g8268 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_111, A2 => lbl2_pxl_n_107, ZN => lbl2_pxl_n_124);
  lbl2_pxl_g8269 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_111, B1 => position_1(10), ZN => lbl2_pxl_n_123);
  lbl2_pxl_g8270 : INR3D0BWP7T port map(A1 => lbl2_pxl_n_88, B1 => lbl2_pxl_n_98, B2 => lbl2_pxl_n_96, ZN => lbl2_pxl_n_122);
  lbl2_pxl_g8271 : AOI211D1BWP7T port map(A1 => lbl2_pxl_n_84, A2 => lbl2_pxl_n_77, B => lbl2_pxl_n_15, C => lbl2_pxl_n_8, ZN => lbl2_pxl_n_121);
  lbl2_pxl_g8272 : OR2D1BWP7T port map(A1 => lbl2_pxl_n_118, A2 => lbl2_pxl_n_8, Z => lbl2_pxl_n_120);
  lbl2_pxl_g8273 : AOI211D1BWP7T port map(A1 => lbl2_pxl_n_79, A2 => lbl2_pxl_n_81, B => lbl2_pxl_n_32, C => lbl2_pxl_n_4, ZN => lbl2_pxl_n_119);
  lbl2_pxl_g8274 : INVD1BWP7T port map(I => lbl2_pxl_n_116, ZN => lbl2_pxl_n_117);
  lbl2_pxl_g8275 : INVD0BWP7T port map(I => lbl2_pxl_n_114, ZN => lbl2_pxl_n_115);
  lbl2_pxl_g8276 : IND2D1BWP7T port map(A1 => player_state_0(0), B1 => lbl2_pxl_n_96, ZN => lbl2_pxl_n_118);
  lbl2_pxl_g8277 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_82, A2 => lbl2_pxl_n_83, B => lbl2_pxl_n_32, ZN => lbl2_pxl_n_116);
  lbl2_pxl_g8278 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_96, B1 => lbl2_pxl_n_98, ZN => lbl2_pxl_n_114);
  lbl2_pxl_g8279 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_78, A2 => lbl2_pxl_n_80, B => lbl2_pxl_n_15, ZN => lbl2_pxl_n_113);
  lbl2_pxl_g8280 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_96, A2 => player_state_0(0), ZN => lbl2_pxl_n_112);
  lbl2_pxl_g8281 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_101, A2 => lbl2_pxl_n_42, ZN => lbl2_pxl_n_111);
  lbl2_pxl_g8282 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_100, B1 => lbl2_data_synced(3), ZN => lbl2_pxl_n_106);
  lbl2_pxl_g8283 : OAI211D1BWP7T port map(A1 => lbl2_pxl_n_42, A2 => lbl2_pxl_n_43, B => lbl2_pxl_n_93, C => lbl2_pxl_n_37, ZN => lbl2_pxl_n_105);
  lbl2_pxl_g8284 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_90, A2 => lbl2_dy_vec(2), B => lbl2_dy_vec(3), ZN => lbl2_pxl_n_110);
  lbl2_pxl_g8285 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_98, A2 => position_1(10), ZN => lbl2_pxl_n_109);
  lbl2_pxl_g8286 : OAI21D0BWP7T port map(A1 => lbl2_pxl_n_89, A2 => lbl2_dy_vec(2), B => lbl2_dy_vec(3), ZN => lbl2_pxl_n_108);
  lbl2_pxl_g8287 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_101, A2 => lbl2_pxl_n_43, ZN => lbl2_pxl_n_107);
  lbl2_pxl_g8288 : INR2D1BWP7T port map(A1 => lbl2_pxl_n_88, B1 => lbl2_pxl_n_91, ZN => lbl2_pxl_n_104);
  lbl2_pxl_g8289 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_92, A2 => lbl2_dx(2), ZN => lbl2_pxl_n_103);
  lbl2_pxl_g8290 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_92, A2 => lbl2_pxl_n_3, ZN => lbl2_pxl_n_102);
  lbl2_pxl_g8291 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_37, B1 => lbl2_pxl_n_90, ZN => lbl2_pxl_n_101);
  lbl2_pxl_g8292 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_65, A2 => lbl2_walls(3), B1 => lbl2_pxl_n_67, B2 => lbl2_walls(2), C => lbl2_pxl_n_86, ZN => lbl2_pxl_n_100);
  lbl2_pxl_g8294 : AOI222D0BWP7T port map(A1 => lbl2_pxl_n_56, A2 => lbl2_pxl_n_55, B1 => lbl2_pxl_n_70, B2 => lbl2_jumps_synced(0), C1 => lbl2_pxl_n_68, C2 => lbl2_jumps_synced(2), ZN => lbl2_pxl_n_95);
  lbl2_pxl_g8295 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_69, A2 => lbl2_jumps_synced(5), B1 => lbl2_pxl_n_71, B2 => lbl2_jumps_synced(7), C => lbl2_pxl_n_76, ZN => lbl2_pxl_n_99);
  lbl2_pxl_g8296 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_93, A2 => lbl2_pxl_n_37, ZN => lbl2_pxl_n_94);
  lbl2_pxl_g8297 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_61, A2 => lbl2_pxl_n_5, B1 => lbl2_pxl_n_62, B2 => direction_1(0), C => lbl2_pxl_n_32, ZN => lbl2_pxl_n_98);
  lbl2_pxl_g8298 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_60, A2 => lbl2_walls(4), B1 => lbl2_pxl_n_59, B2 => lbl2_walls(6), C => lbl2_pxl_n_85, ZN => lbl2_pxl_n_97);
  lbl2_pxl_g8299 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_61, A2 => lbl2_pxl_n_10, B1 => lbl2_pxl_n_62, B2 => direction_0(0), C => lbl2_pxl_n_15, ZN => lbl2_pxl_n_96);
  lbl2_pxl_g8300 : INVD0BWP7T port map(I => lbl2_pxl_n_90, ZN => lbl2_pxl_n_89);
  lbl2_pxl_g8301 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_75, A2 => lbl2_pxl_n_38, ZN => lbl2_pxl_n_93);
  lbl2_pxl_g8302 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_69, A2 => lbl2_jumps_synced(1), B1 => lbl2_pxl_n_71, B2 => lbl2_jumps_synced(3), ZN => lbl2_pxl_n_87);
  lbl2_pxl_g8303 : AO22D0BWP7T port map(A1 => lbl2_pxl_n_63, A2 => lbl2_walls(1), B1 => lbl2_walls(0), B2 => lbl2_pxl_n_66, Z => lbl2_pxl_n_86);
  lbl2_pxl_g8304 : AO22D0BWP7T port map(A1 => lbl2_pxl_n_57, A2 => lbl2_walls(5), B1 => lbl2_walls(7), B2 => lbl2_pxl_n_58, Z => lbl2_pxl_n_85);
  lbl2_pxl_g8305 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_37, B1 => lbl2_pxl_n_75, ZN => lbl2_pxl_n_92);
  lbl2_pxl_g8306 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_49, A2 => lbl2_borders_synced(4), B1 => lbl2_pxl_n_51, B2 => lbl2_borders_synced(7), C => lbl2_pxl_n_73, ZN => lbl2_pxl_n_91);
  lbl2_pxl_g8307 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_74, A2 => lbl2_pxl_n_53, ZN => lbl2_pxl_n_90);
  lbl2_pxl_g8308 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_49, A2 => lbl2_borders_synced(0), B1 => lbl2_pxl_n_51, B2 => lbl2_borders_synced(3), C => lbl2_pxl_n_72, ZN => lbl2_pxl_n_88);
  lbl2_pxl_g8309 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_59, A2 => lbl2_pxl_n_20, B1 => lbl2_pxl_n_58, B2 => lbl2_pxl_n_26, ZN => lbl2_pxl_n_84);
  lbl2_pxl_g8310 : AOI33D1BWP7T port map(A1 => lbl2_pxl_n_66, A2 => lbl2_pxl_n_5, A3 => direction_1(1), B1 => lbl2_pxl_n_63, B2 => direction_1(0), B3 => direction_1(1), ZN => lbl2_pxl_n_83);
  lbl2_pxl_g8311 : MAOI22D0BWP7T port map(A1 => lbl2_pxl_n_67, A2 => lbl2_pxl_n_25, B1 => lbl2_pxl_n_64, B2 => lbl2_pxl_n_29, ZN => lbl2_pxl_n_82);
  lbl2_pxl_g8312 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_57, A2 => lbl2_pxl_n_17, B1 => lbl2_pxl_n_58, B2 => lbl2_pxl_n_28, ZN => lbl2_pxl_n_81);
  lbl2_pxl_g8313 : MAOI22D0BWP7T port map(A1 => lbl2_pxl_n_63, A2 => lbl2_pxl_n_24, B1 => lbl2_pxl_n_64, B2 => lbl2_pxl_n_27, ZN => lbl2_pxl_n_80);
  lbl2_pxl_g8314 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_60, A2 => lbl2_pxl_n_31, B1 => lbl2_pxl_n_59, B2 => lbl2_pxl_n_25, ZN => lbl2_pxl_n_79);
  lbl2_pxl_g8315 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_67, A2 => lbl2_pxl_n_20, B1 => lbl2_pxl_n_66, B2 => lbl2_pxl_n_19, ZN => lbl2_pxl_n_78);
  lbl2_pxl_g8316 : AOI33D1BWP7T port map(A1 => lbl2_pxl_n_60, A2 => lbl2_pxl_n_10, A3 => direction_0(1), B1 => lbl2_pxl_n_57, B2 => direction_0(0), B3 => direction_0(1), ZN => lbl2_pxl_n_77);
  lbl2_pxl_g8317 : AO22D0BWP7T port map(A1 => lbl2_pxl_n_70, A2 => lbl2_jumps_synced(4), B1 => lbl2_jumps_synced(6), B2 => lbl2_pxl_n_68, Z => lbl2_pxl_n_76);
  lbl2_pxl_g8318 : INVD0BWP7T port map(I => lbl2_pxl_n_74, ZN => lbl2_pxl_n_75);
  lbl2_pxl_g8319 : MAOI222D1BWP7T port map(A => lbl2_pxl_n_46, B => lbl2_pxl_n_35, C => lbl2_pxl_n_34, ZN => lbl2_pxl_n_74);
  lbl2_pxl_g8320 : AO22D0BWP7T port map(A1 => lbl2_pxl_n_50, A2 => lbl2_borders_synced(5), B1 => lbl2_borders_synced(6), B2 => lbl2_pxl_n_52, Z => lbl2_pxl_n_73);
  lbl2_pxl_g8321 : AO22D0BWP7T port map(A1 => lbl2_pxl_n_50, A2 => lbl2_borders_synced(1), B1 => lbl2_borders_synced(2), B2 => lbl2_pxl_n_52, Z => lbl2_pxl_n_72);
  lbl2_pxl_g8322 : INVD0BWP7T port map(I => lbl2_pxl_n_64, ZN => lbl2_pxl_n_65);
  lbl2_pxl_g8323 : AO21D0BWP7T port map(A1 => lbl2_pxl_n_39, A2 => lbl2_dy_vec(1), B => lbl2_pxl_n_51, Z => lbl2_pxl_n_71);
  lbl2_pxl_g8324 : AO21D0BWP7T port map(A1 => lbl2_pxl_n_41, A2 => lbl2_dx(1), B => lbl2_pxl_n_49, Z => lbl2_pxl_n_70);
  lbl2_pxl_g8325 : AO21D0BWP7T port map(A1 => lbl2_pxl_n_40, A2 => lbl2_dy_vec(1), B => lbl2_pxl_n_50, Z => lbl2_pxl_n_69);
  lbl2_pxl_g8326 : AO21D0BWP7T port map(A1 => lbl2_pxl_n_44, A2 => lbl2_dx(1), B => lbl2_pxl_n_52, Z => lbl2_pxl_n_68);
  lbl2_pxl_g8327 : IAO21D0BWP7T port map(A1 => lbl2_dy_vec(3), A2 => lbl2_dy_vec(2), B => lbl2_pxl_n_38, ZN => lbl2_pxl_n_67);
  lbl2_pxl_g8328 : AOI21D0BWP7T port map(A1 => lbl2_dy_vec(3), A2 => lbl2_dy_vec(2), B => lbl2_pxl_n_38, ZN => lbl2_pxl_n_66);
  lbl2_pxl_g8329 : OAI21D0BWP7T port map(A1 => lbl2_dx(3), A2 => lbl2_dx(2), B => lbl2_pxl_n_37, ZN => lbl2_pxl_n_64);
  lbl2_pxl_g8330 : OA21D0BWP7T port map(A1 => lbl2_pxl_n_6, A2 => lbl2_pxl_n_3, B => lbl2_pxl_n_37, Z => lbl2_pxl_n_63);
  lbl2_pxl_g8331 : OAI33D1BWP7T port map(A1 => lbl2_dx(0), A2 => lbl2_pxl_n_6, A3 => lbl2_pxl_n_12, B1 => lbl2_pxl_n_9, B2 => lbl2_dx(3), B3 => lbl2_pxl_n_14, ZN => lbl2_pxl_n_56);
  lbl2_pxl_g8332 : OAI33D1BWP7T port map(A1 => lbl2_dy_vec(0), A2 => lbl2_pxl_n_7, A3 => lbl2_pxl_n_13, B1 => lbl2_pxl_n_11, B2 => lbl2_dy_vec(3), B3 => lbl2_pxl_n_22, ZN => lbl2_pxl_n_55);
  lbl2_pxl_g8333 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_42, A2 => position_1(10), B1 => lbl2_pxl_n_43, B2 => position_0(10), ZN => lbl2_pxl_n_54);
  lbl2_pxl_g8334 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_45, A2 => lbl2_pxl_n_37, ZN => lbl2_pxl_n_62);
  lbl2_pxl_g8335 : OR3XD1BWP7T port map(A1 => lbl2_pxl_n_44, A2 => lbl2_pxl_n_41, A3 => lbl2_pxl_n_38, Z => lbl2_pxl_n_61);
  lbl2_pxl_g8336 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_13, A2 => lbl2_dy_vec(3), B => lbl2_pxl_n_47, ZN => lbl2_pxl_n_60);
  lbl2_pxl_g8337 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_22, A2 => lbl2_pxl_n_7, B => lbl2_pxl_n_47, ZN => lbl2_pxl_n_59);
  lbl2_pxl_g8338 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_14, A2 => lbl2_pxl_n_6, B => lbl2_pxl_n_48, ZN => lbl2_pxl_n_58);
  lbl2_pxl_g8339 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_12, A2 => lbl2_dx(3), B => lbl2_pxl_n_48, ZN => lbl2_pxl_n_57);
  lbl2_pxl_g8340 : INVD0BWP7T port map(I => lbl2_pxl_n_38, ZN => lbl2_pxl_n_53);
  lbl2_pxl_g8341 : AN2D1BWP7T port map(A1 => lbl2_pxl_n_44, A2 => lbl2_dy_vec(0), Z => lbl2_pxl_n_52);
  lbl2_pxl_g8342 : AN2D1BWP7T port map(A1 => lbl2_pxl_n_39, A2 => lbl2_dx(0), Z => lbl2_pxl_n_51);
  lbl2_pxl_g8343 : AN2D1BWP7T port map(A1 => lbl2_pxl_n_40, A2 => lbl2_pxl_n_9, Z => lbl2_pxl_n_50);
  lbl2_pxl_g8344 : AN2D1BWP7T port map(A1 => lbl2_pxl_n_41, A2 => lbl2_pxl_n_11, Z => lbl2_pxl_n_49);
  lbl2_pxl_g8345 : OAI221D0BWP7T port map(A1 => lbl2_dx(2), A2 => lbl2_dx(0), B1 => lbl2_pxl_n_9, B2 => lbl2_pxl_n_3, C => lbl2_pxl_n_36, ZN => lbl2_pxl_n_46);
  lbl2_pxl_g8346 : NR2D0BWP7T port map(A1 => lbl2_pxl_n_40, A2 => lbl2_pxl_n_39, ZN => lbl2_pxl_n_45);
  lbl2_pxl_g8347 : OA22D0BWP7T port map(A1 => lbl2_pxl_n_13, A2 => lbl2_pxl_n_7, B1 => lbl2_dy_vec(3), B2 => lbl2_pxl_n_22, Z => lbl2_pxl_n_48);
  lbl2_pxl_g8348 : OA22D0BWP7T port map(A1 => lbl2_pxl_n_12, A2 => lbl2_pxl_n_6, B1 => lbl2_dx(3), B2 => lbl2_pxl_n_14, Z => lbl2_pxl_n_47);
  lbl2_pxl_g8349 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_22, A2 => lbl2_pxl_n_7, ZN => lbl2_pxl_n_44);
  lbl2_pxl_g8350 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_21, A2 => player_state_0(0), ZN => lbl2_pxl_n_43);
  lbl2_pxl_g8351 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_33, A2 => player_state_1(0), ZN => lbl2_pxl_n_42);
  lbl2_pxl_g8352 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_13, A2 => lbl2_dy_vec(3), ZN => lbl2_pxl_n_41);
  lbl2_pxl_g8355 : MAOI22D0BWP7T port map(A1 => lbl2_dy_vec(2), A2 => lbl2_dy_vec(0), B1 => lbl2_dy_vec(2), B2 => lbl2_dy_vec(0), ZN => lbl2_pxl_n_36);
  lbl2_pxl_g8356 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_12, A2 => lbl2_pxl_n_14, ZN => lbl2_pxl_n_35);
  lbl2_pxl_g8357 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_13, A2 => lbl2_pxl_n_22, ZN => lbl2_pxl_n_34);
  lbl2_pxl_g8358 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_12, A2 => lbl2_dx(3), ZN => lbl2_pxl_n_40);
  lbl2_pxl_g8359 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_14, A2 => lbl2_pxl_n_6, ZN => lbl2_pxl_n_39);
  lbl2_pxl_g8360 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_3, A2 => lbl2_dx(3), B1 => lbl2_pxl_n_6, B2 => lbl2_dx(2), ZN => lbl2_pxl_n_38);
  lbl2_pxl_g8361 : MOAI22D0BWP7T port map(A1 => lbl2_pxl_n_7, A2 => lbl2_dy_vec(2), B1 => lbl2_pxl_n_7, B2 => lbl2_dy_vec(2), ZN => lbl2_pxl_n_37);
  lbl2_pxl_g8363 : INVD0BWP7T port map(I => lbl2_pxl_n_30, ZN => lbl2_pxl_n_31);
  lbl2_pxl_g8364 : CKND1BWP7T port map(I => lbl2_pxl_n_28, ZN => lbl2_pxl_n_29);
  lbl2_pxl_g8365 : CKND1BWP7T port map(I => lbl2_pxl_n_26, ZN => lbl2_pxl_n_27);
  lbl2_pxl_g8366 : INVD0BWP7T port map(I => lbl2_pxl_n_23, ZN => lbl2_pxl_n_24);
  lbl2_pxl_g8367 : IND2D1BWP7T port map(A1 => player_state_1(1), B1 => lbl2_n_189, ZN => lbl2_pxl_n_33);
  lbl2_pxl_g8368 : ND2D1BWP7T port map(A1 => lbl2_n_189, A2 => player_state_1(1), ZN => lbl2_pxl_n_32);
  lbl2_pxl_g8369 : CKND2D1BWP7T port map(A1 => lbl2_pxl_n_5, A2 => direction_1(1), ZN => lbl2_pxl_n_30);
  lbl2_pxl_g8370 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_5, A2 => direction_1(1), ZN => lbl2_pxl_n_28);
  lbl2_pxl_g8371 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_10, A2 => direction_0(1), ZN => lbl2_pxl_n_26);
  lbl2_pxl_g8372 : NR2D0BWP7T port map(A1 => direction_1(1), A2 => direction_1(0), ZN => lbl2_pxl_n_25);
  lbl2_pxl_g8373 : CKND2D1BWP7T port map(A1 => direction_0(1), A2 => direction_0(0), ZN => lbl2_pxl_n_23);
  lbl2_pxl_g8374 : CKND2D1BWP7T port map(A1 => lbl2_dy_vec(2), A2 => lbl2_dy_vec(1), ZN => lbl2_pxl_n_22);
  lbl2_pxl_g8376 : INVD0BWP7T port map(I => lbl2_pxl_n_18, ZN => lbl2_pxl_n_19);
  lbl2_pxl_g8377 : INVD0BWP7T port map(I => lbl2_pxl_n_16, ZN => lbl2_pxl_n_17);
  lbl2_pxl_g8378 : IND2D1BWP7T port map(A1 => player_state_0(1), B1 => lbl2_n_190, ZN => lbl2_pxl_n_21);
  lbl2_pxl_g8379 : NR2D0BWP7T port map(A1 => direction_0(1), A2 => direction_0(0), ZN => lbl2_pxl_n_20);
  lbl2_pxl_g8380 : CKND2D1BWP7T port map(A1 => lbl2_pxl_n_10, A2 => direction_0(1), ZN => lbl2_pxl_n_18);
  lbl2_pxl_g8381 : CKND2D1BWP7T port map(A1 => direction_1(1), A2 => direction_1(0), ZN => lbl2_pxl_n_16);
  lbl2_pxl_g8382 : ND2D1BWP7T port map(A1 => lbl2_n_190, A2 => player_state_0(1), ZN => lbl2_pxl_n_15);
  lbl2_pxl_g8383 : ND2D1BWP7T port map(A1 => lbl2_dx(1), A2 => lbl2_dx(2), ZN => lbl2_pxl_n_14);
  lbl2_pxl_g8384 : OR2D1BWP7T port map(A1 => lbl2_dy_vec(1), A2 => lbl2_dy_vec(2), Z => lbl2_pxl_n_13);
  lbl2_pxl_g8385 : IND2D1BWP7T port map(A1 => lbl2_dx(1), B1 => lbl2_pxl_n_3, ZN => lbl2_pxl_n_12);
  lbl2_pxl_g8386 : INVD0BWP7T port map(I => lbl2_dy_vec(0), ZN => lbl2_pxl_n_11);
  lbl2_pxl_g8387 : INVD1BWP7T port map(I => direction_0(0), ZN => lbl2_pxl_n_10);
  lbl2_pxl_g8388 : INVD1BWP7T port map(I => lbl2_dx(0), ZN => lbl2_pxl_n_9);
  lbl2_pxl_g8389 : INVD1BWP7T port map(I => position_0(10), ZN => lbl2_pxl_n_8);
  lbl2_pxl_g8390 : INVD1BWP7T port map(I => lbl2_dy_vec(3), ZN => lbl2_pxl_n_7);
  lbl2_pxl_g8391 : INVD1BWP7T port map(I => lbl2_dx(3), ZN => lbl2_pxl_n_6);
  lbl2_pxl_g8392 : INVD1BWP7T port map(I => direction_1(0), ZN => lbl2_pxl_n_5);
  lbl2_pxl_g8393 : INVD0BWP7T port map(I => position_1(10), ZN => lbl2_pxl_n_4);
  lbl2_pxl_g8394 : INVD1BWP7T port map(I => lbl2_dx(2), ZN => lbl2_pxl_n_3);
  lbl2_pxl_g2 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_97, B1 => lbl2_pxl_n_172, B2 => lbl2_data_synced(7), ZN => lbl2_pxl_n_2);
  lbl2_pxl_g8395 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_33, B1 => player_state_1(0), ZN => lbl2_pxl_n_1);
  lbl2_pxl_g8396 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_21, B1 => player_state_0(0), ZN => lbl2_pxl_n_0);
  lbl2_sdb_g8069 : OR2D1BWP7T port map(A1 => lbl2_sidebar_color(3), A2 => lbl2_sdb_n_167, Z => lbl2_sidebar_color(2));
  lbl2_sdb_g8070 : OR2D1BWP7T port map(A1 => lbl2_sidebar_color(1), A2 => lbl2_sdb_n_167, Z => lbl2_sidebar_color(0));
  lbl2_sdb_g8071 : AN2D0BWP7T port map(A1 => lbl2_sdb_n_179, A2 => lbl2_h_count(9), Z => lbl2_sidebar_color(3));
  lbl2_sdb_g8072 : INR2D1BWP7T port map(A1 => lbl2_sdb_n_179, B1 => lbl2_h_count(9), ZN => lbl2_sidebar_color(1));
  lbl2_sdb_g8073 : OAI211D1BWP7T port map(A1 => lbl2_v_count(7), A2 => lbl2_sdb_n_178, B => lbl2_sdb_n_176, C => lbl2_sdb_n_160, ZN => lbl2_sdb_n_179);
  lbl2_sdb_g8074 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_177, A2 => lbl2_v_count(5), ZN => lbl2_sdb_n_178);
  lbl2_sdb_g8075 : NR4D0BWP7T port map(A1 => lbl2_sdb_n_175, A2 => game_state(2), A3 => lbl2_v_count(8), A4 => lbl2_v_count(6), ZN => lbl2_sdb_n_177);
  lbl2_sdb_g8076 : NR4D0BWP7T port map(A1 => lbl2_sdb_n_173, A2 => lbl2_sdb_n_169, A3 => lbl2_sdb_n_170, A4 => lbl2_sdb_n_151, ZN => lbl2_sdb_n_176);
  lbl2_sdb_g8077 : AOI31D0BWP7T port map(A1 => lbl2_sdb_n_163, A2 => lbl2_sdb_n_31, A3 => game_state(1), B => lbl2_sdb_n_174, ZN => lbl2_sdb_n_175);
  lbl2_sdb_g8078 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_172, A2 => lbl2_sdb_n_161, B => lbl2_sdb_n_79, ZN => lbl2_sdb_n_174);
  lbl2_sdb_g8079 : OAI32D1BWP7T port map(A1 => lbl2_sdb_n_16, A2 => lbl2_sdb_n_79, A3 => lbl2_sdb_n_171, B1 => lbl2_sdb_n_33, B2 => lbl2_sdb_n_124, ZN => lbl2_sdb_n_173);
  lbl2_sdb_g8080 : IND3D1BWP7T port map(A1 => lbl2_sdb_n_31, B1 => game_state(1), B2 => lbl2_sdb_n_168, ZN => lbl2_sdb_n_172);
  lbl2_sdb_g8081 : OAI211D1BWP7T port map(A1 => lbl2_sdb_n_139, A2 => lbl2_sdb_n_164, B => lbl2_sdb_n_32, C => lbl2_sdb_n_43, ZN => lbl2_sdb_n_171);
  lbl2_sdb_g8082 : NR3D0BWP7T port map(A1 => lbl2_sdb_n_166, A2 => lbl2_sdb_n_63, A3 => lbl2_h_count(9), ZN => lbl2_sdb_n_170);
  lbl2_sdb_g8083 : OAI32D1BWP7T port map(A1 => lbl2_v_count(5), A2 => lbl2_sdb_n_16, A3 => lbl2_sdb_n_122, B1 => lbl2_sdb_n_6, B2 => lbl2_sdb_n_165, ZN => lbl2_sdb_n_169);
  lbl2_sdb_g8084 : OAI221D0BWP7T port map(A1 => lbl2_sdb_n_142, A2 => lbl2_sdb_n_29, B1 => lbl2_sdb_n_36, B2 => lbl2_sdb_n_93, C => lbl2_sdb_n_162, ZN => lbl2_sdb_n_168);
  lbl2_sdb_g8085 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_165, A2 => lbl2_n_152, ZN => lbl2_sdb_n_167);
  lbl2_sdb_g8086 : OA32D1BWP7T port map(A1 => lbl2_sdb_n_29, A2 => lbl2_sdb_n_79, A3 => lbl2_sdb_n_0, B1 => lbl2_sdb_n_79, B2 => lbl2_sdb_n_149, Z => lbl2_sdb_n_166);
  lbl2_sdb_g8087 : AOI221D0BWP7T port map(A1 => lbl2_sdb_n_155, A2 => lbl2_sdb_n_29, B1 => lbl2_sdb_n_130, B2 => lbl2_sdb_n_108, C => lbl2_sdb_n_146, ZN => lbl2_sdb_n_164);
  lbl2_sdb_g8088 : IND4D0BWP7T port map(A1 => lbl2_sdb_n_158, B1 => lbl2_v_count(6), B2 => lbl2_v_count(5), B3 => lbl2_v_count(7), ZN => lbl2_sdb_n_165);
  lbl2_sdb_g8089 : AOI211D1BWP7T port map(A1 => lbl2_sdb_n_55, A2 => lbl2_n_151, B => lbl2_sdb_n_159, C => lbl2_sdb_n_65, ZN => lbl2_sdb_n_163);
  lbl2_sdb_g8090 : AOI211XD0BWP7T port map(A1 => lbl2_sdb_n_157, A2 => lbl2_sdb_n_29, B => lbl2_sdb_n_152, C => lbl2_sdb_n_140, ZN => lbl2_sdb_n_162);
  lbl2_sdb_g8091 : OAI31D0BWP7T port map(A1 => lbl2_sdb_n_120, A2 => lbl2_sdb_n_143, A3 => lbl2_sdb_n_153, B => lbl2_sdb_n_28, ZN => lbl2_sdb_n_161);
  lbl2_sdb_g8092 : IND3D1BWP7T port map(A1 => lbl2_sdb_n_63, B1 => lbl2_h_count(9), B2 => lbl2_sdb_n_156, ZN => lbl2_sdb_n_160);
  lbl2_sdb_g8094 : AOI211XD0BWP7T port map(A1 => lbl2_sdb_n_148, A2 => lbl2_h_count(2), B => lbl2_sdb_n_141, C => lbl2_sdb_n_138, ZN => lbl2_sdb_n_159);
  lbl2_sdb_g8095 : IND4D0BWP7T port map(A1 => lbl2_v_count(8), B1 => game_state(2), B2 => lbl2_sdb_n_28, B3 => lbl2_sdb_n_131, ZN => lbl2_sdb_n_158);
  lbl2_sdb_g8096 : OAI221D0BWP7T port map(A1 => lbl2_sdb_n_136, A2 => lbl2_sdb_n_81, B1 => lbl2_sdb_n_84, B2 => lbl2_sdb_n_108, C => lbl2_sdb_n_144, ZN => lbl2_sdb_n_157);
  lbl2_sdb_g8097 : OAI221D0BWP7T port map(A1 => lbl2_sdb_n_52, A2 => lbl2_sdb_n_82, B1 => lbl2_sdb_n_77, B2 => lbl2_sdb_n_60, C => lbl2_sdb_n_150, ZN => lbl2_sdb_n_156);
  lbl2_sdb_g8098 : OA211D0BWP7T port map(A1 => lbl2_sdb_n_77, A2 => lbl2_sdb_n_108, B => lbl2_sdb_n_154, C => lbl2_sdb_n_94, Z => lbl2_sdb_n_155);
  lbl2_sdb_g8099 : OA221D0BWP7T port map(A1 => lbl2_sdb_n_109, A2 => lbl2_sdb_n_62, B1 => lbl2_sdb_n_24, B2 => lbl2_sdb_n_93, C => lbl2_sdb_n_145, Z => lbl2_sdb_n_154);
  lbl2_sdb_g8100 : OAI211D1BWP7T port map(A1 => lbl2_sdb_n_94, A2 => lbl2_sdb_n_128, B => lbl2_sdb_n_135, C => lbl2_sdb_n_119, ZN => lbl2_sdb_n_153);
  lbl2_sdb_g8101 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_137, A2 => lbl2_sdb_n_92, B => lbl2_sdb_n_57, ZN => lbl2_sdb_n_152);
  lbl2_sdb_g8102 : OAI33D1BWP7T port map(A1 => lbl2_sdb_n_15, A2 => lbl2_n_151, A3 => lbl2_sdb_n_126, B1 => lbl2_sdb_n_2, B2 => lbl2_sdb_n_17, B3 => lbl2_sdb_n_117, ZN => lbl2_sdb_n_151);
  lbl2_sdb_g8103 : AOI211XD0BWP7T port map(A1 => lbl2_sdb_n_125, A2 => lbl2_sdb_n_29, B => lbl2_sdb_n_98, C => lbl2_sdb_n_96, ZN => lbl2_sdb_n_150);
  lbl2_sdb_g8104 : MAOI22D0BWP7T port map(A1 => lbl2_sdb_n_134, A2 => lbl2_sdb_n_13, B1 => lbl2_sdb_n_127, B2 => lbl2_sdb_n_82, ZN => lbl2_sdb_n_149);
  lbl2_sdb_g8105 : OAI32D1BWP7T port map(A1 => lbl2_v_count(4), A2 => lbl2_sdb_n_30, A3 => lbl2_sdb_n_89, B1 => lbl2_sdb_n_75, B2 => lbl2_sdb_n_133, ZN => lbl2_sdb_n_148);
  lbl2_sdb_g8106 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_121, A2 => lbl2_sdb_n_110, B => lbl2_sdb_n_44, ZN => lbl2_sdb_n_147);
  lbl2_sdb_g8107 : OA211D0BWP7T port map(A1 => lbl2_sdb_n_92, A2 => lbl2_sdb_n_112, B => lbl2_sdb_n_93, C => lbl2_sdb_n_50, Z => lbl2_sdb_n_146);
  lbl2_sdb_g8108 : AOI33D1BWP7T port map(A1 => lbl2_sdb_n_114, A2 => lbl2_sdb_n_90, A3 => lbl2_v_count(2), B1 => lbl2_sdb_n_113, B2 => lbl2_sdb_n_84, B3 => lbl2_sdb_n_13, ZN => lbl2_sdb_n_145);
  lbl2_sdb_g8110 : MOAI22D0BWP7T port map(A1 => lbl2_sdb_n_127, A2 => lbl2_sdb_n_90, B1 => lbl2_sdb_n_129, B2 => lbl2_sdb_n_29, ZN => lbl2_sdb_n_143);
  lbl2_sdb_g8111 : OA22D0BWP7T port map(A1 => lbl2_sdb_n_127, A2 => lbl2_sdb_n_62, B1 => lbl2_sdb_n_19, B2 => lbl2_sdb_n_92, Z => lbl2_sdb_n_142);
  lbl2_sdb_g8112 : AOI33D1BWP7T port map(A1 => lbl2_sdb_n_113, A2 => lbl2_sdb_n_70, A3 => lbl2_v_count(2), B1 => lbl2_sdb_n_77, B2 => lbl2_sdb_n_13, B3 => lbl2_sdb_n_7, ZN => lbl2_sdb_n_144);
  lbl2_sdb_g8113 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_123, A2 => lbl2_h_count(2), ZN => lbl2_sdb_n_141);
  lbl2_sdb_g8114 : NR2D0BWP7T port map(A1 => lbl2_sdb_n_128, A2 => lbl2_sdb_n_93, ZN => lbl2_sdb_n_140);
  lbl2_sdb_g8115 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_109, A2 => lbl2_sdb_n_111, B => lbl2_sdb_n_92, ZN => lbl2_sdb_n_139);
  lbl2_sdb_g8116 : OA221D0BWP7T port map(A1 => lbl2_sdb_n_105, A2 => lbl2_sdb_n_83, B1 => lbl2_sdb_n_18, B2 => lbl2_sdb_n_30, C => lbl2_sdb_n_118, Z => lbl2_sdb_n_138);
  lbl2_sdb_g8117 : OA31D1BWP7T port map(A1 => FE_DBTN0_lbl2_v_count_2, A2 => lbl2_sdb_n_90, A3 => lbl2_sdb_n_103, B => lbl2_sdb_n_110, Z => lbl2_sdb_n_137);
  lbl2_sdb_g8118 : AOI31D0BWP7T port map(A1 => lbl2_sdb_n_103, A2 => lbl2_sdb_n_84, A3 => lbl2_sdb_n_35, B => lbl2_sdb_n_114, ZN => lbl2_sdb_n_136);
  lbl2_sdb_g8119 : AO211D0BWP7T port map(A1 => lbl2_sdb_n_84, A2 => lbl2_sdb_n_29, B => lbl2_sdb_n_109, C => lbl2_sdb_n_77, Z => lbl2_sdb_n_135);
  lbl2_sdb_g8120 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_92, A2 => lbl2_sdb_n_90, B => lbl2_sdb_n_128, ZN => lbl2_sdb_n_134);
  lbl2_sdb_g8121 : AOI222D0BWP7T port map(A1 => lbl2_sdb_n_105, A2 => lbl2_sdb_n_30, B1 => lbl2_sdb_n_100, B2 => lbl2_sdb_n_7, C1 => lbl2_sdb_n_89, C2 => lbl2_sdb_n_20, ZN => lbl2_sdb_n_133);
  lbl2_sdb_g8122 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_109, A2 => lbl2_sdb_n_112, B => lbl2_sdb_n_62, ZN => lbl2_sdb_n_132);
  lbl2_sdb_g8123 : OAI221D0BWP7T port map(A1 => lbl2_sdb_n_106, A2 => lbl2_sdb_n_50, B1 => lbl2_sdb_n_77, B2 => lbl2_sdb_n_69, C => lbl2_sdb_n_107, ZN => lbl2_sdb_n_131);
  lbl2_sdb_g8124 : OAI32D1BWP7T port map(A1 => FE_DBTN0_lbl2_v_count_2, A2 => lbl2_sdb_n_29, A3 => lbl2_sdb_n_91, B1 => lbl2_sdb_n_29, B2 => lbl2_sdb_n_113, ZN => lbl2_sdb_n_130);
  lbl2_sdb_g8125 : IAO21D0BWP7T port map(A1 => lbl2_sdb_n_71, A2 => lbl2_n_154, B => lbl2_sdb_n_116, ZN => lbl2_sdb_n_126);
  lbl2_sdb_g8126 : OAI211D1BWP7T port map(A1 => lbl2_v_count(3), A2 => lbl2_sdb_n_87, B => lbl2_sdb_n_85, C => lbl2_sdb_n_48, ZN => lbl2_sdb_n_125);
  lbl2_sdb_g8127 : IAO21D0BWP7T port map(A1 => lbl2_sdb_n_74, A2 => lbl2_n_154, B => lbl2_sdb_n_115, ZN => lbl2_sdb_n_124);
  lbl2_sdb_g8128 : INR2D1BWP7T port map(A1 => lbl2_sdb_n_114, B1 => lbl2_sdb_n_90, ZN => lbl2_sdb_n_129);
  lbl2_sdb_g8129 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_113, A2 => lbl2_sdb_n_29, ZN => lbl2_sdb_n_128);
  lbl2_sdb_g8130 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_114, A2 => FE_DBTN0_lbl2_v_count_2, ZN => lbl2_sdb_n_127);
  lbl2_sdb_g8131 : AOI22D0BWP7T port map(A1 => lbl2_sdb_n_95, A2 => lbl2_sdb_n_88, B1 => lbl2_sdb_n_97, B2 => lbl2_sdb_n_49, ZN => lbl2_sdb_n_123);
  lbl2_sdb_g8132 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_73, A2 => lbl2_n_154, B => lbl2_sdb_n_115, ZN => lbl2_sdb_n_122);
  lbl2_sdb_g8133 : OAI21D0BWP7T port map(A1 => lbl2_sdb_n_104, A2 => lbl2_sdb_n_37, B => lbl2_sdb_n_84, ZN => lbl2_sdb_n_121);
  lbl2_sdb_g8134 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_90, A2 => lbl2_sdb_n_82, B => lbl2_sdb_n_108, ZN => lbl2_sdb_n_120);
  lbl2_sdb_g8135 : IOA21D1BWP7T port map(A1 => lbl2_sdb_n_80, A2 => lbl2_sdb_n_81, B => lbl2_sdb_n_113, ZN => lbl2_sdb_n_119);
  lbl2_sdb_g8136 : MAOI22D0BWP7T port map(A1 => lbl2_sdb_n_102, A2 => lbl2_sdb_n_83, B1 => lbl2_sdb_n_75, B2 => lbl2_sdb_n_13, ZN => lbl2_sdb_n_118);
  lbl2_sdb_g8137 : AOI31D0BWP7T port map(A1 => lbl2_sdb_n_68, A2 => lbl2_n_154, A3 => lbl2_n_153, B => lbl2_sdb_n_116, ZN => lbl2_sdb_n_117);
  lbl2_sdb_g8138 : INVD0BWP7T port map(I => lbl2_sdb_n_113, ZN => lbl2_sdb_n_112);
  lbl2_sdb_g8139 : CKND2D0BWP7T port map(A1 => lbl2_sdb_n_104, A2 => lbl2_sdb_n_37, ZN => lbl2_sdb_n_111);
  lbl2_sdb_g8140 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_99, A2 => lbl2_sdb_n_56, ZN => lbl2_sdb_n_116);
  lbl2_sdb_g8141 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_54, A2 => lbl2_sdb_n_99, ZN => lbl2_sdb_n_115);
  lbl2_sdb_g8142 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_103, A2 => lbl2_v_count(4), ZN => lbl2_sdb_n_114);
  lbl2_sdb_g8143 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_104, A2 => lbl2_v_count(4), ZN => lbl2_sdb_n_113);
  lbl2_sdb_g8144 : OA33D0BWP7T port map(A1 => lbl2_sdb_n_44, A2 => lbl2_sdb_n_80, A3 => lbl2_sdb_n_38, B1 => lbl2_sdb_n_29, B2 => lbl2_sdb_n_81, B3 => lbl2_sdb_n_21, Z => lbl2_sdb_n_107);
  lbl2_sdb_g8145 : OA221D0BWP7T port map(A1 => lbl2_sdb_n_64, A2 => lbl2_n_149, B1 => lbl2_sdb_n_24, B2 => lbl2_sdb_n_17, C => lbl2_sdb_n_101, Z => lbl2_sdb_n_106);
  lbl2_sdb_g8146 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_103, A2 => lbl2_sdb_n_70, ZN => lbl2_sdb_n_110);
  lbl2_sdb_g8147 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_103, A2 => lbl2_sdb_n_20, ZN => lbl2_sdb_n_109);
  lbl2_sdb_g8148 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_104, A2 => lbl2_sdb_n_20, ZN => lbl2_sdb_n_108);
  lbl2_sdb_g8149 : INVD1BWP7T port map(I => lbl2_sdb_n_104, ZN => lbl2_sdb_n_103);
  lbl2_sdb_g8150 : ND2D0BWP7T port map(A1 => lbl2_sdb_n_88, A2 => lbl2_sdb_n_20, ZN => lbl2_sdb_n_102);
  lbl2_sdb_g8151 : IAO21D0BWP7T port map(A1 => lbl2_sdb_n_39, A2 => lbl2_sdb_n_15, B => lbl2_sdb_n_86, ZN => lbl2_sdb_n_101);
  lbl2_sdb_g8152 : NR2D0BWP7T port map(A1 => lbl2_sdb_n_89, A2 => lbl2_sdb_n_27, ZN => lbl2_sdb_n_100);
  lbl2_sdb_g8153 : NR2D0BWP7T port map(A1 => lbl2_sdb_n_88, A2 => lbl2_v_count(4), ZN => lbl2_sdb_n_105);
  lbl2_sdb_g8154 : IOA21D1BWP7T port map(A1 => lbl2_sdb_n_67, A2 => lbl2_n_150, B => lbl2_sdb_n_66, ZN => lbl2_sdb_n_104);
  lbl2_sdb_g8155 : NR3D0BWP7T port map(A1 => lbl2_sdb_n_21, A2 => lbl2_sdb_n_80, A3 => lbl2_v_count(2), ZN => lbl2_sdb_n_98);
  lbl2_sdb_g8156 : AOI211XD0BWP7T port map(A1 => lbl2_sdb_n_19, A2 => lbl2_v_count(4), B => lbl2_sdb_n_88, C => lbl2_sdb_n_76, ZN => lbl2_sdb_n_97);
  lbl2_sdb_g8157 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_81, A2 => lbl2_sdb_n_57, B => lbl2_sdb_n_38, ZN => lbl2_sdb_n_96);
  lbl2_sdb_g8158 : OAI32D1BWP7T port map(A1 => FE_DBTN2_lbl2_h_count_3, A2 => lbl2_v_count(4), A3 => lbl2_sdb_n_76, B1 => lbl2_sdb_n_36, B2 => lbl2_sdb_n_75, ZN => lbl2_sdb_n_95);
  lbl2_sdb_g8159 : AOI222D0BWP7T port map(A1 => lbl2_sdb_n_42, A2 => lbl2_sdb_n_61, B1 => lbl2_sdb_n_41, B2 => lbl2_sdb_n_30, C1 => lbl2_sdb_n_78, C2 => lbl2_sdb_n_34, ZN => lbl2_sdb_n_99);
  lbl2_sdb_g8160 : INVD0BWP7T port map(I => lbl2_sdb_n_92, ZN => lbl2_sdb_n_91);
  lbl2_sdb_g8161 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_70, A2 => lbl2_sdb_n_20, ZN => lbl2_sdb_n_94);
  lbl2_sdb_g8162 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_84, A2 => lbl2_sdb_n_77, ZN => lbl2_sdb_n_93);
  lbl2_sdb_g8163 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_70, A2 => lbl2_sdb_n_77, ZN => lbl2_sdb_n_92);
  lbl2_sdb_g8164 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_84, A2 => lbl2_sdb_n_62, ZN => lbl2_sdb_n_90);
  lbl2_sdb_g8165 : INVD1BWP7T port map(I => lbl2_sdb_n_89, ZN => lbl2_sdb_n_88);
  lbl2_sdb_g8166 : AO21D0BWP7T port map(A1 => lbl2_sdb_n_15, A2 => lbl2_sdb_n_77, B => lbl2_sdb_n_40, Z => lbl2_sdb_n_87);
  lbl2_sdb_g8167 : IAO21D0BWP7T port map(A1 => lbl2_sdb_n_15, A2 => lbl2_sdb_n_62, B => lbl2_sdb_n_40, ZN => lbl2_sdb_n_86);
  lbl2_sdb_g8168 : AOI22D0BWP7T port map(A1 => lbl2_sdb_n_51, A2 => lbl2_sdb_n_62, B1 => lbl2_sdb_n_46, B2 => lbl2_v_count(2), ZN => lbl2_sdb_n_85);
  lbl2_sdb_g8169 : OAI21D0BWP7T port map(A1 => lbl2_sdb_n_72, A2 => lbl2_sdb_n_10, B => lbl2_sdb_n_55, ZN => lbl2_sdb_n_89);
  lbl2_sdb_g8170 : INVD1BWP7T port map(I => lbl2_sdb_n_70, ZN => lbl2_sdb_n_84);
  lbl2_sdb_g8171 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_76, A2 => lbl2_sdb_n_49, ZN => lbl2_sdb_n_83);
  lbl2_sdb_g8172 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_77, A2 => lbl2_sdb_n_29, ZN => lbl2_sdb_n_82);
  lbl2_sdb_g8173 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_62, A2 => lbl2_sdb_n_20, ZN => lbl2_sdb_n_81);
  lbl2_sdb_g8174 : MOAI22D0BWP7T port map(A1 => lbl2_sdb_n_12, A2 => FE_DBTN1_lbl2_h_count_1, B1 => lbl2_sdb_n_14, B2 => FE_DBTN2_lbl2_h_count_3, ZN => lbl2_sdb_n_78);
  lbl2_sdb_g8175 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_62, A2 => lbl2_sdb_n_50, ZN => lbl2_sdb_n_80);
  lbl2_sdb_g8176 : MOAI22D0BWP7T port map(A1 => lbl2_sdb_n_66, A2 => lbl2_n_151, B1 => lbl2_sdb_n_66, B2 => lbl2_n_151, ZN => lbl2_sdb_n_79);
  lbl2_sdb_g8177 : INVD1BWP7T port map(I => lbl2_sdb_n_62, ZN => lbl2_sdb_n_77);
  lbl2_sdb_g8178 : INVD1BWP7T port map(I => lbl2_sdb_n_76, ZN => lbl2_sdb_n_75);
  lbl2_sdb_g8179 : CKND1BWP7T port map(I => lbl2_sdb_n_73, ZN => lbl2_sdb_n_74);
  lbl2_sdb_g8180 : HA1D0BWP7T port map(A => lbl2_sdb_n_12, B => lbl2_sdb_n_2, CO => lbl2_sdb_n_72, S => lbl2_sdb_n_76);
  lbl2_sdb_g8181 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_68, A2 => lbl2_n_153, ZN => lbl2_sdb_n_71);
  lbl2_sdb_g8182 : NR3D0BWP7T port map(A1 => lbl2_sdb_n_54, A2 => lbl2_sdb_n_58, A3 => lbl2_n_153, ZN => lbl2_sdb_n_73);
  lbl2_sdb_g8183 : IAO21D0BWP7T port map(A1 => lbl2_sdb_n_39, A2 => lbl2_sdb_n_2, B => lbl2_sdb_n_59, ZN => lbl2_sdb_n_69);
  lbl2_sdb_g8184 : OAI21D0BWP7T port map(A1 => lbl2_sdb_n_2, A2 => lbl2_sdb_n_53, B => lbl2_sdb_n_67, ZN => lbl2_sdb_n_70);
  lbl2_sdb_g8185 : NR2D0BWP7T port map(A1 => lbl2_sdb_n_56, A2 => lbl2_sdb_n_58, ZN => lbl2_sdb_n_68);
  lbl2_sdb_g8186 : NR2XD0BWP7T port map(A1 => lbl2_sdb_n_55, A2 => lbl2_n_151, ZN => lbl2_sdb_n_65);
  lbl2_sdb_g8187 : OAI21D0BWP7T port map(A1 => lbl2_sdb_n_46, A2 => lbl2_sdb_n_45, B => lbl2_sdb_n_9, ZN => lbl2_sdb_n_64);
  lbl2_sdb_g8188 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_2, A2 => lbl2_sdb_n_53, ZN => lbl2_sdb_n_67);
  lbl2_sdb_g8189 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_26, A2 => lbl2_sdb_n_53, ZN => lbl2_sdb_n_66);
  lbl2_sdb_g8190 : OAI32D1BWP7T port map(A1 => lbl2_h_count(2), A2 => lbl2_h_count(3), A3 => FE_DBTN1_lbl2_h_count_1, B1 => lbl2_h_count(1), B2 => lbl2_sdb_n_12, ZN => lbl2_sdb_n_61);
  lbl2_sdb_g8191 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_45, A2 => lbl2_sdb_n_2, B => lbl2_sdb_n_47, ZN => lbl2_sdb_n_60);
  lbl2_sdb_g8192 : AO33D0BWP7T port map(A1 => lbl2_sdb_n_8, A2 => lbl2_sdb_n_2, A3 => lbl2_sdb_n_37, B1 => lbl2_sdb_n_22, B2 => lbl2_sdb_n_10, B3 => FE_DBTN0_lbl2_v_count_2, Z => lbl2_sdb_n_59);
  lbl2_sdb_g8193 : IND3D1BWP7T port map(A1 => lbl2_sdb_n_43, B1 => lbl2_sdb_n_5, B2 => lbl2_sdb_n_32, ZN => lbl2_sdb_n_63);
  lbl2_sdb_g8194 : MOAI22D1BWP7T port map(A1 => lbl2_sdb_n_14, A2 => lbl2_h_count(3), B1 => lbl2_sdb_n_14, B2 => lbl2_h_count(3), ZN => lbl2_sdb_n_62);
  lbl2_sdb_g8195 : NR2XD0BWP7T port map(A1 => lbl2_sdb_n_34, A2 => lbl2_sdb_n_30, ZN => lbl2_sdb_n_58);
  lbl2_sdb_g8196 : IND2D1BWP7T port map(A1 => lbl2_sdb_n_24, B1 => lbl2_sdb_n_29, ZN => lbl2_sdb_n_57);
  lbl2_sdb_g8197 : IND3D1BWP7T port map(A1 => lbl2_sdb_n_33, B1 => lbl2_v_count(7), B2 => lbl2_v_count(4), ZN => lbl2_sdb_n_56);
  lbl2_sdb_g8198 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_26, A2 => lbl2_sdb_n_12, ZN => lbl2_sdb_n_55);
  lbl2_sdb_g8199 : AOI33D1BWP7T port map(A1 => lbl2_sdb_n_22, A2 => lbl2_sdb_n_2, A3 => lbl2_sdb_n_20, B1 => lbl2_sdb_n_26, B2 => lbl2_sdb_n_23, B3 => lbl2_v_count(2), ZN => lbl2_sdb_n_52);
  lbl2_sdb_g8200 : AO21D0BWP7T port map(A1 => lbl2_sdb_n_22, A2 => lbl2_sdb_n_25, B => lbl2_sdb_n_45, Z => lbl2_sdb_n_51);
  lbl2_sdb_g8201 : IND4D0BWP7T port map(A1 => lbl2_sdb_n_17, B1 => lbl2_v_count(7), B2 => lbl2_sdb_n_7, B3 => lbl2_sdb_n_2, ZN => lbl2_sdb_n_54);
  lbl2_sdb_g8202 : OA21D0BWP7T port map(A1 => FE_DBTN1_lbl2_h_count_1, A2 => FE_DBTN2_lbl2_h_count_3, B => lbl2_sdb_n_12, Z => lbl2_sdb_n_53);
  lbl2_sdb_g8203 : INVD0BWP7T port map(I => lbl2_sdb_n_29, ZN => lbl2_sdb_n_50);
  lbl2_sdb_g8204 : INVD0BWP7T port map(I => lbl2_sdb_n_30, ZN => lbl2_sdb_n_49);
  lbl2_sdb_g8205 : CKND1BWP7T port map(I => lbl2_sdb_n_47, ZN => lbl2_sdb_n_48);
  lbl2_sdb_g8206 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_39, A2 => lbl2_sdb_n_10, ZN => lbl2_sdb_n_47);
  lbl2_sdb_g8207 : NR2D0BWP7T port map(A1 => lbl2_sdb_n_38, A2 => lbl2_v_count(4), ZN => lbl2_sdb_n_46);
  lbl2_sdb_g8208 : NR2D1BWP7T port map(A1 => lbl2_n_151, A2 => lbl2_sdb_n_36, ZN => lbl2_sdb_n_45);
  lbl2_sdb_g8209 : MOAI22D0BWP7T port map(A1 => lbl2_sdb_n_27, A2 => lbl2_v_count(1), B1 => lbl2_sdb_n_20, B2 => lbl2_v_count(1), ZN => lbl2_sdb_n_42);
  lbl2_sdb_g8210 : MUX2ND0BWP7T port map(I0 => lbl2_sdb_n_19, I1 => lbl2_sdb_n_27, S => lbl2_v_count(1), ZN => lbl2_sdb_n_41);
  lbl2_sdb_g8211 : NR2XD0BWP7T port map(A1 => lbl2_sdb_n_35, A2 => lbl2_sdb_n_23, ZN => lbl2_sdb_n_44);
  lbl2_sdb_g8212 : OA21D0BWP7T port map(A1 => lbl2_sdb_n_16, A2 => lbl2_sdb_n_11, B => lbl2_sdb_n_5, Z => lbl2_sdb_n_43);
  lbl2_sdb_g8213 : CKND1BWP7T port map(I => lbl2_sdb_n_36, ZN => lbl2_sdb_n_35);
  lbl2_sdb_g8214 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_22, A2 => lbl2_v_count(2), ZN => lbl2_sdb_n_40);
  lbl2_sdb_g8215 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_8, A2 => lbl2_sdb_n_20, ZN => lbl2_sdb_n_39);
  lbl2_sdb_g8216 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_26, A2 => lbl2_n_151, ZN => lbl2_sdb_n_38);
  lbl2_sdb_g8217 : NR2D0BWP7T port map(A1 => lbl2_sdb_n_24, A2 => lbl2_v_count(2), ZN => lbl2_sdb_n_37);
  lbl2_sdb_g8218 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_20, A2 => lbl2_v_count(4), ZN => lbl2_sdb_n_36);
  lbl2_sdb_g8219 : OR2D1BWP7T port map(A1 => lbl2_sdb_n_18, A2 => lbl2_sdb_n_13, Z => lbl2_sdb_n_34);
  lbl2_sdb_g8220 : IND3D0BWP7T port map(A1 => lbl2_v_count(6), B1 => lbl2_v_count(8), B2 => lbl2_v_count(5), ZN => lbl2_sdb_n_33);
  lbl2_sdb_g8221 : NR3D0BWP7T port map(A1 => game_state(0), A2 => game_state(1), A3 => game_state(2), ZN => lbl2_sdb_n_32);
  lbl2_sdb_g8222 : MOAI22D0BWP7T port map(A1 => game_state(0), A2 => lbl2_h_count(9), B1 => game_state(0), B2 => lbl2_h_count(9), ZN => lbl2_sdb_n_31);
  lbl2_sdb_g8223 : MOAI22D0BWP7T port map(A1 => FE_DBTN2_lbl2_h_count_3, A2 => lbl2_h_count(2), B1 => FE_DBTN2_lbl2_h_count_3, B2 => lbl2_h_count(2), ZN => lbl2_sdb_n_30);
  lbl2_sdb_g8224 : AOI21D1BWP7T port map(A1 => lbl2_h_count(1), A2 => lbl2_h_count(2), B => lbl2_sdb_n_14, ZN => lbl2_sdb_n_29);
  lbl2_sdb_g8225 : INVD0BWP7T port map(I => lbl2_sdb_n_26, ZN => lbl2_sdb_n_25);
  lbl2_sdb_g8226 : INVD0BWP7T port map(I => lbl2_sdb_n_24, ZN => lbl2_sdb_n_23);
  lbl2_sdb_g8227 : INVD0BWP7T port map(I => lbl2_sdb_n_22, ZN => lbl2_sdb_n_21);
  lbl2_sdb_g8228 : INVD0BWP7T port map(I => lbl2_sdb_n_20, ZN => lbl2_sdb_n_19);
  lbl2_sdb_g8229 : INR2D1BWP7T port map(A1 => game_state(0), B1 => game_state(1), ZN => lbl2_sdb_n_28);
  lbl2_sdb_g8230 : ND2D1BWP7T port map(A1 => lbl2_v_count(2), A2 => lbl2_v_count(3), ZN => lbl2_sdb_n_27);
  lbl2_sdb_g8231 : NR2XD0BWP7T port map(A1 => lbl2_n_150, A2 => lbl2_n_149, ZN => lbl2_sdb_n_26);
  lbl2_sdb_g8232 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_7, A2 => lbl2_v_count(3), ZN => lbl2_sdb_n_24);
  lbl2_sdb_g8233 : NR2D1BWP7T port map(A1 => lbl2_n_151, A2 => lbl2_v_count(4), ZN => lbl2_sdb_n_22);
  lbl2_sdb_g8234 : NR2XD0BWP7T port map(A1 => lbl2_v_count(2), A2 => lbl2_v_count(3), ZN => lbl2_sdb_n_20);
  lbl2_sdb_g8235 : NR2D0BWP7T port map(A1 => lbl2_sdb_n_9, A2 => lbl2_v_count(2), ZN => lbl2_sdb_n_18);
  lbl2_sdb_g8236 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_8, A2 => lbl2_n_150, ZN => lbl2_sdb_n_17);
  lbl2_sdb_g8237 : CKND2D1BWP7T port map(A1 => lbl2_v_count(8), A2 => lbl2_v_count(6), ZN => lbl2_sdb_n_16);
  lbl2_sdb_g8238 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_10, A2 => lbl2_n_149, ZN => lbl2_sdb_n_15);
  lbl2_sdb_g8239 : NR2D1BWP7T port map(A1 => lbl2_h_count(1), A2 => lbl2_h_count(2), ZN => lbl2_sdb_n_14);
  lbl2_sdb_g8240 : NR2D1BWP7T port map(A1 => FE_DBTN0_lbl2_v_count_2, A2 => lbl2_v_count(3), ZN => lbl2_sdb_n_13);
  lbl2_sdb_g8241 : ND2D1BWP7T port map(A1 => lbl2_h_count(2), A2 => lbl2_h_count(3), ZN => lbl2_sdb_n_12);
  lbl2_sdb_g8242 : INVD0BWP7T port map(I => lbl2_v_count(5), ZN => lbl2_sdb_n_11);
  lbl2_sdb_g8243 : INVD1BWP7T port map(I => lbl2_n_150, ZN => lbl2_sdb_n_10);
  lbl2_sdb_g8244 : INVD0BWP7T port map(I => lbl2_v_count(3), ZN => lbl2_sdb_n_9);
  lbl2_sdb_g8245 : INVD1BWP7T port map(I => lbl2_n_151, ZN => lbl2_sdb_n_8);
  lbl2_sdb_g8246 : INVD1BWP7T port map(I => lbl2_v_count(4), ZN => lbl2_sdb_n_7);
  lbl2_sdb_g8247 : CKND1BWP7T port map(I => lbl2_n_152, ZN => lbl2_sdb_n_6);
  lbl2_sdb_g8248 : INVD0BWP7T port map(I => lbl2_v_count(7), ZN => lbl2_sdb_n_5);
  lbl2_sdb_g8251 : INVD1BWP7T port map(I => lbl2_n_149, ZN => lbl2_sdb_n_2);
  lbl2_sdb_g2 : INR4D0BWP7T port map(A1 => lbl2_sdb_n_144, B1 => lbl2_sdb_n_147, B2 => lbl2_sdb_n_132, B3 => lbl2_sdb_n_129, ZN => lbl2_sdb_n_0);
  lbl0_g14543 : IND4D0BWP7T port map(A1 => lbl0_n_422, B1 => lbl0_n_245, B2 => lbl0_n_362, B3 => lbl0_n_408, ZN => lbl0_n_416);
  lbl0_g14544 : IND4D0BWP7T port map(A1 => lbl0_n_422, B1 => lbl0_n_248, B2 => lbl0_n_361, B3 => lbl0_n_408, ZN => lbl0_n_415);
  lbl0_g14545 : AOI31D0BWP7T port map(A1 => lbl0_n_406, A2 => lbl0_n_221, A3 => lbl0_n_199, B => lbl0_n_407, ZN => lbl0_n_408);
  lbl0_g14546 : IND3D1BWP7T port map(A1 => lbl0_n_407, B1 => lbl0_n_248, B2 => lbl0_n_264, ZN => lbl0_n_420);
  lbl0_g14547 : IND3D1BWP7T port map(A1 => lbl0_n_407, B1 => lbl0_n_245, B2 => lbl0_n_263, ZN => lbl0_n_421);
  lbl0_g14548 : AOI211D1BWP7T port map(A1 => lbl0_n_402, A2 => position_0(9), B => lbl0_n_405, C => lbl0_n_403, ZN => lbl0_n_407);
  lbl0_g14549 : NR4D0BWP7T port map(A1 => lbl0_n_404, A2 => lbl0_n_397, A3 => lbl0_n_391, A4 => lbl0_n_379, ZN => lbl0_n_406);
  lbl0_g14550 : IND4D0BWP7T port map(A1 => lbl0_n_399, B1 => lbl0_n_221, B2 => lbl0_n_394, B3 => lbl0_n_401, ZN => lbl0_n_405);
  lbl0_g14551 : OAI21D0BWP7T port map(A1 => lbl0_n_402, A2 => lbl0_n_279, B => lbl0_n_220, ZN => lbl0_d_position_1(9));
  lbl0_g14552 : MOAI22D0BWP7T port map(A1 => lbl0_n_402, A2 => lbl0_n_400, B1 => lbl0_n_402, B2 => lbl0_n_400, ZN => lbl0_n_404);
  lbl0_g14553 : NR2XD0BWP7T port map(A1 => lbl0_n_402, A2 => position_0(9), ZN => lbl0_n_403);
  lbl0_g14554 : OAI221D0BWP7T port map(A1 => lbl0_n_396, A2 => lbl0_n_316, B1 => lbl0_n_318, B2 => lbl0_n_398, C => lbl0_n_390, ZN => address(9));
  lbl0_g14555 : AN2D0BWP7T port map(A1 => lbl0_n_400, A2 => lbl0_n_281, Z => lbl0_n_414);
  lbl0_g14556 : MAOI22D0BWP7T port map(A1 => lbl0_next_direction_1(0), A2 => position_1(9), B1 => lbl0_n_398, B2 => lbl0_next_direction_1(0), ZN => lbl0_n_402);
  lbl0_g14557 : AOI211XD0BWP7T port map(A1 => lbl0_n_388, A2 => position_0(8), B => lbl0_n_395, C => lbl0_n_369, ZN => lbl0_n_401);
  lbl0_g14558 : MOAI22D0BWP7T port map(A1 => lbl0_n_396, A2 => lbl0_next_direction_0(0), B1 => lbl0_next_direction_0(0), B2 => position_0(9), ZN => lbl0_n_400);
  lbl0_g14559 : OAI21D0BWP7T port map(A1 => lbl0_n_388, A2 => lbl0_n_279, B => lbl0_n_168, ZN => lbl0_d_position_1(8));
  lbl0_g14560 : OAI211D1BWP7T port map(A1 => position_0(8), A2 => lbl0_n_388, B => lbl0_n_135, C => lbl0_n_196, ZN => lbl0_n_399);
  lbl0_g14561 : MOAI22D0BWP7T port map(A1 => lbl0_n_388, A2 => lbl0_n_385, B1 => lbl0_n_388, B2 => lbl0_n_385, ZN => lbl0_n_397);
  lbl0_g14562 : MAOI22D0BWP7T port map(A1 => lbl0_n_389, A2 => position_1(9), B1 => lbl0_n_389, B2 => position_1(9), ZN => lbl0_n_398);
  lbl0_g14563 : OAI221D0BWP7T port map(A1 => lbl0_n_350, A2 => lbl0_n_316, B1 => lbl0_n_318, B2 => lbl0_n_359, C => lbl0_n_387, ZN => address(7));
  lbl0_g14564 : OAI221D0BWP7T port map(A1 => lbl0_n_373, A2 => lbl0_n_316, B1 => lbl0_n_318, B2 => lbl0_n_377, C => lbl0_n_386, ZN => address(8));
  lbl0_g14565 : ND2D1BWP7T port map(A1 => lbl0_n_393, A2 => lbl0_n_346, ZN => address(6));
  lbl0_g14566 : OAI221D0BWP7T port map(A1 => lbl0_n_316, A2 => position_0(5), B1 => position_1(5), B2 => lbl0_n_318, C => lbl0_n_392, ZN => address(5));
  lbl0_g14567 : MOAI22D0BWP7T port map(A1 => lbl0_n_385, A2 => lbl0_n_158, B1 => lbl0_n_385, B2 => lbl0_n_158, ZN => lbl0_n_395);
  lbl0_g14568 : AO21D0BWP7T port map(A1 => lbl0_n_385, A2 => lbl0_n_281, B => lbl0_n_215, Z => lbl0_d_position_0(8));
  lbl0_g14569 : NR4D0BWP7T port map(A1 => lbl0_n_380, A2 => lbl0_n_383, A3 => lbl0_n_376, A4 => lbl0_n_259, ZN => lbl0_n_394);
  lbl0_g14570 : MAOI22D0BWP7T port map(A1 => lbl0_n_384, A2 => position_0(9), B1 => lbl0_n_384, B2 => position_0(9), ZN => lbl0_n_396);
  lbl0_g14571 : AOI22D0BWP7T port map(A1 => lbl0_n_381, A2 => position_1(6), B1 => lbl0_n_336, B2 => position_0(6), ZN => lbl0_n_393);
  lbl0_g14572 : AOI22D0BWP7T port map(A1 => lbl0_n_381, A2 => position_1(5), B1 => lbl0_n_336, B2 => position_0(5), ZN => lbl0_n_392);
  lbl0_g14573 : ND4D0BWP7T port map(A1 => lbl0_n_382, A2 => lbl0_n_355, A3 => lbl0_n_367, A4 => lbl0_n_366, ZN => lbl0_n_391);
  lbl0_g14574 : AOI22D0BWP7T port map(A1 => lbl0_n_381, A2 => position_1(9), B1 => lbl0_n_336, B2 => position_0(9), ZN => lbl0_n_390);
  lbl0_g14575 : AOI22D0BWP7T port map(A1 => lbl0_n_381, A2 => position_1(7), B1 => lbl0_n_336, B2 => position_0(7), ZN => lbl0_n_387);
  lbl0_g14576 : AOI22D0BWP7T port map(A1 => lbl0_n_381, A2 => position_1(8), B1 => lbl0_n_336, B2 => position_0(8), ZN => lbl0_n_386);
  lbl0_g14577 : MAOI22D0BWP7T port map(A1 => lbl0_n_378, A2 => lbl0_n_167, B1 => lbl0_n_378, B2 => lbl0_n_167, ZN => lbl0_n_389);
  lbl0_g14578 : MAOI22D0BWP7T port map(A1 => lbl0_next_direction_1(0), A2 => position_1(8), B1 => lbl0_n_377, B2 => lbl0_next_direction_1(0), ZN => lbl0_n_388);
  lbl0_g14579 : OAI21D0BWP7T port map(A1 => lbl0_n_371, A2 => lbl0_n_279, B => lbl0_n_168, ZN => lbl0_d_position_1(7));
  lbl0_g14580 : MOAI22D0BWP7T port map(A1 => lbl0_n_373, A2 => lbl0_next_direction_0(0), B1 => lbl0_next_direction_0(0), B2 => position_0(8), ZN => lbl0_n_385);
  lbl0_g14581 : MOAI22D0BWP7T port map(A1 => lbl0_n_371, A2 => position_0(7), B1 => lbl0_n_371, B2 => position_0(7), ZN => lbl0_n_383);
  lbl0_g14582 : MAOI22D0BWP7T port map(A1 => lbl0_n_371, A2 => lbl0_n_368, B1 => lbl0_n_371, B2 => lbl0_n_368, ZN => lbl0_n_382);
  lbl0_g14583 : MAOI22D0BWP7T port map(A1 => lbl0_n_372, A2 => lbl0_n_181, B1 => lbl0_n_372, B2 => lbl0_n_181, ZN => lbl0_n_384);
  lbl0_g14584 : OAI221D0BWP7T port map(A1 => lbl0_n_348, A2 => position_0(4), B1 => position_0(5), B2 => lbl0_n_204, C => lbl0_n_375, ZN => lbl0_n_380);
  lbl0_g14585 : ND4D0BWP7T port map(A1 => lbl0_n_356, A2 => lbl0_n_354, A3 => lbl0_n_353, A4 => lbl0_n_258, ZN => lbl0_n_379);
  lbl0_g14586 : INR2XD0BWP7T port map(A1 => lbl0_n_374, B1 => lbl0_state(4), ZN => lbl0_n_381);
  lbl0_g14587 : AO21D0BWP7T port map(A1 => lbl0_n_368, A2 => lbl0_n_281, B => lbl0_n_215, Z => lbl0_d_position_0(7));
  lbl0_g14588 : AOI22D0BWP7T port map(A1 => lbl0_n_352, A2 => lbl0_n_167, B1 => lbl0_n_312, B2 => position_1(8), ZN => lbl0_n_378);
  lbl0_g14589 : AOI22D0BWP7T port map(A1 => lbl0_n_360, A2 => lbl0_n_167, B1 => lbl0_n_342, B2 => lbl0_n_166, ZN => lbl0_n_377);
  lbl0_g14590 : OAI221D0BWP7T port map(A1 => lbl0_n_338, A2 => position_0(2), B1 => position_0(1), B2 => lbl0_n_296, C => lbl0_n_370, ZN => lbl0_n_376);
  lbl0_g14591 : AOI221D0BWP7T port map(A1 => lbl0_n_348, A2 => position_0(4), B1 => lbl0_n_204, B2 => position_0(5), C => lbl0_n_357, ZN => lbl0_n_375);
  lbl0_g14592 : NR4D0BWP7T port map(A1 => lbl0_n_351, A2 => lbl0_n_336, A3 => lbl0_n_317, A4 => lbl0_n_319, ZN => lbl0_n_374);
  lbl0_g14593 : OAI221D0BWP7T port map(A1 => lbl0_n_349, A2 => lbl0_n_299, B1 => lbl0_n_302, B2 => lbl0_n_348, C => lbl0_n_335, ZN => address(4));
  lbl0_g14594 : MAOI22D0BWP7T port map(A1 => lbl0_n_324, A2 => lbl0_n_181, B1 => lbl0_n_365, B2 => lbl0_n_181, ZN => lbl0_n_373);
  lbl0_g14595 : OAI22D0BWP7T port map(A1 => lbl0_n_364, A2 => lbl0_n_181, B1 => lbl0_n_297, B2 => lbl0_n_159, ZN => lbl0_n_372);
  lbl0_g14596 : MAOI22D0BWP7T port map(A1 => lbl0_next_direction_1(0), A2 => position_1(7), B1 => lbl0_n_359, B2 => lbl0_next_direction_1(0), ZN => lbl0_n_371);
  lbl0_g14597 : OAI221D0BWP7T port map(A1 => lbl0_n_331, A2 => lbl0_n_299, B1 => lbl0_n_302, B2 => lbl0_n_330, C => lbl0_n_329, ZN => address(3));
  lbl0_g14598 : AOI221D0BWP7T port map(A1 => lbl0_n_338, A2 => position_0(2), B1 => lbl0_n_296, B2 => position_0(1), C => lbl0_n_358, ZN => lbl0_n_370);
  lbl0_g14599 : OAI221D0BWP7T port map(A1 => lbl0_n_294, A2 => position_1(1), B1 => position_1(5), B2 => lbl0_n_202, C => lbl0_n_363, ZN => lbl0_n_369);
  lbl0_g14600 : OAI221D0BWP7T port map(A1 => lbl0_n_340, A2 => lbl0_n_299, B1 => lbl0_n_302, B2 => lbl0_n_338, C => lbl0_n_328, ZN => address(2));
  lbl0_g14601 : AOI22D0BWP7T port map(A1 => lbl0_n_349, A2 => lbl0_n_347, B1 => lbl0_n_204, B2 => lbl0_n_201, ZN => lbl0_n_367);
  lbl0_g14602 : MAOI22D0BWP7T port map(A1 => lbl0_n_202, A2 => lbl0_n_203, B1 => lbl0_n_349, B2 => lbl0_n_347, ZN => lbl0_n_366);
  lbl0_g14603 : OAI22D0BWP7T port map(A1 => lbl0_n_348, A2 => lbl0_n_279, B1 => lbl0_n_168, B2 => start_position_0(3), ZN => lbl0_d_position_1(4));
  lbl0_g14604 : MOAI22D0BWP7T port map(A1 => lbl0_n_350, A2 => lbl0_next_direction_0(0), B1 => lbl0_next_direction_0(0), B2 => position_0(7), ZN => lbl0_n_368);
  lbl0_g14605 : HA1D0BWP7T port map(A => lbl0_n_159, B => lbl0_n_315, CO => lbl0_n_364, S => lbl0_n_365);
  lbl0_g14606 : NR2D1BWP7T port map(A1 => lbl0_n_349, A2 => lbl0_n_280, ZN => lbl0_n_412);
  lbl0_g14607 : AOI221D0BWP7T port map(A1 => lbl0_n_294, A2 => position_1(1), B1 => lbl0_n_202, B2 => position_1(5), C => lbl0_n_344, ZN => lbl0_n_363);
  lbl0_g14608 : ND3D0BWP7T port map(A1 => lbl0_n_325, A2 => lbl0_n_427, A3 => lbl0_n_241, ZN => lbl0_n_362);
  lbl0_g14609 : ND3D0BWP7T port map(A1 => lbl0_n_323, A2 => lbl0_n_427, A3 => lbl0_n_227, ZN => lbl0_n_361);
  lbl0_g14610 : OAI21D0BWP7T port map(A1 => lbl0_n_340, A2 => lbl0_n_280, B => lbl0_n_220, ZN => lbl0_d_position_0(2));
  lbl0_g14611 : OAI222D0BWP7T port map(A1 => lbl0_n_321, A2 => lbl0_n_155, B1 => lbl0_n_262, B2 => lbl0_n_143, C1 => lbl0_n_261, C2 => lbl0_n_306, ZN => write_memory(4));
  lbl0_g14612 : OAI21D0BWP7T port map(A1 => lbl0_n_339, A2 => lbl0_n_279, B => lbl0_n_216, ZN => lbl0_d_position_1(6));
  lbl0_g14613 : OAI21D0BWP7T port map(A1 => lbl0_n_341, A2 => lbl0_n_158, B => lbl0_n_352, ZN => lbl0_n_360);
  lbl0_g14614 : OAI21D0BWP7T port map(A1 => lbl0_n_338, A2 => lbl0_n_279, B => lbl0_n_168, ZN => lbl0_d_position_1(2));
  lbl0_g14615 : OAI21D0BWP7T port map(A1 => lbl0_n_306, A2 => lbl0_n_208, B => lbl0_n_343, ZN => write_memory(6));
  lbl0_g14616 : OAI21D0BWP7T port map(A1 => lbl0_n_307, A2 => lbl0_n_208, B => lbl0_n_345, ZN => write_memory(2));
  lbl0_g14617 : MOAI22D0BWP7T port map(A1 => lbl0_n_330, A2 => lbl0_n_279, B1 => lbl0_n_505, B2 => start_position_1(3), ZN => lbl0_d_position_1(3));
  lbl0_g14618 : MOAI22D0BWP7T port map(A1 => lbl0_n_331, A2 => lbl0_n_280, B1 => lbl0_n_505, B2 => start_position_0(3), ZN => lbl0_d_position_0(3));
  lbl0_g14619 : MOAI22D0BWP7T port map(A1 => lbl0_n_330, A2 => position_0(3), B1 => lbl0_n_330, B2 => position_0(3), ZN => lbl0_n_358);
  lbl0_g14620 : MOAI22D0BWP7T port map(A1 => lbl0_n_339, A2 => position_0(6), B1 => lbl0_n_339, B2 => position_0(6), ZN => lbl0_n_357);
  lbl0_g14621 : XNR2D1BWP7T port map(A1 => lbl0_n_330, A2 => lbl0_n_331, ZN => lbl0_n_356);
  lbl0_g14622 : XNR2D1BWP7T port map(A1 => lbl0_n_339, A2 => lbl0_n_311, ZN => lbl0_n_355);
  lbl0_g14623 : MAOI22D0BWP7T port map(A1 => lbl0_n_294, A2 => lbl0_n_295, B1 => lbl0_n_337, B2 => lbl0_n_340, ZN => lbl0_n_354);
  lbl0_g14624 : AOI22D0BWP7T port map(A1 => lbl0_n_337, A2 => lbl0_n_340, B1 => lbl0_n_296, B2 => lbl0_n_293, ZN => lbl0_n_353);
  lbl0_g14625 : MAOI22D0BWP7T port map(A1 => lbl0_n_332, A2 => position_1(7), B1 => lbl0_n_332, B2 => position_1(7), ZN => lbl0_n_359);
  lbl0_g14626 : OAI222D0BWP7T port map(A1 => lbl0_n_321, A2 => lbl0_n_163, B1 => lbl0_n_240, B2 => lbl0_n_306, C1 => lbl0_n_243, C2 => lbl0_n_143, ZN => write_memory(5));
  lbl0_g14627 : OAI221D0BWP7T port map(A1 => lbl0_n_294, A2 => lbl0_n_299, B1 => lbl0_n_302, B2 => lbl0_n_296, C => lbl0_n_326, ZN => address(1));
  lbl0_g14628 : IND4D0BWP7T port map(A1 => lbl0_n_426, B1 => lbl0_n_419, B2 => lbl0_n_282, B3 => lbl0_n_292, ZN => lbl0_n_351);
  lbl0_g14629 : OAI21D0BWP7T port map(A1 => lbl0_n_321, A2 => lbl0_n_164, B => lbl0_n_143, ZN => write_memory(7));
  lbl0_g14630 : OAI221D0BWP7T port map(A1 => lbl0_n_299, A2 => lbl0_n_205, B1 => lbl0_n_200, B2 => lbl0_n_302, C => lbl0_n_327, ZN => address(0));
  lbl0_g14631 : AO21D0BWP7T port map(A1 => lbl0_n_322, A2 => lbl0_read_data_reg(3), B => lbl0_n_305, Z => write_memory(3));
  lbl0_g14632 : OAI221D0BWP7T port map(A1 => lbl0_n_307, A2 => lbl0_n_261, B1 => lbl0_n_262, B2 => lbl0_n_304, C => lbl0_n_334, ZN => write_memory(0));
  lbl0_g14633 : OAI21D0BWP7T port map(A1 => lbl0_n_311, A2 => lbl0_n_280, B => lbl0_n_216, ZN => lbl0_d_position_0(6));
  lbl0_g14634 : ND2D1BWP7T port map(A1 => lbl0_n_341, A2 => lbl0_n_158, ZN => lbl0_n_352);
  lbl0_g14635 : INVD0BWP7T port map(I => lbl0_n_348, ZN => lbl0_n_347);
  lbl0_g14636 : AOI22D0BWP7T port map(A1 => lbl0_n_319, A2 => lbl0_n_276, B1 => lbl0_n_317, B2 => lbl0_n_287, ZN => lbl0_n_346);
  lbl0_g14637 : AOI22D0BWP7T port map(A1 => lbl0_n_322, A2 => lbl0_read_data_reg(2), B1 => lbl0_n_305, B2 => lbl0_n_207, ZN => lbl0_n_345);
  lbl0_g14638 : OAI221D0BWP7T port map(A1 => lbl0_n_307, A2 => lbl0_n_240, B1 => lbl0_n_243, B2 => lbl0_n_304, C => lbl0_n_333, ZN => write_memory(1));
  lbl0_g14639 : MOAI22D0BWP7T port map(A1 => lbl0_n_311, A2 => position_1(6), B1 => lbl0_n_311, B2 => position_1(6), ZN => lbl0_n_344);
  lbl0_g14640 : MAOI22D0BWP7T port map(A1 => lbl0_n_320, A2 => lbl0_read_data_reg(6), B1 => lbl0_n_143, B2 => lbl0_n_249, ZN => lbl0_n_343);
  lbl0_g14641 : MOAI22D0BWP7T port map(A1 => lbl0_n_312, A2 => lbl0_n_158, B1 => lbl0_n_312, B2 => lbl0_n_158, ZN => lbl0_n_342);
  lbl0_g14642 : MAOI22D0BWP7T port map(A1 => lbl0_n_313, A2 => position_0(7), B1 => lbl0_n_313, B2 => position_0(7), ZN => lbl0_n_350);
  lbl0_g14643 : MAOI22D0BWP7T port map(A1 => lbl0_n_137, A2 => position_0(4), B1 => lbl0_n_137, B2 => position_0(4), ZN => lbl0_n_349);
  lbl0_g14644 : MAOI22D0BWP7T port map(A1 => lbl0_n_314, A2 => position_1(4), B1 => lbl0_n_314, B2 => position_1(4), ZN => lbl0_n_348);
  lbl0_g14645 : INVD0BWP7T port map(I => lbl0_n_338, ZN => lbl0_n_337);
  lbl0_g14646 : AOI22D0BWP7T port map(A1 => lbl0_n_301, A2 => position_0(4), B1 => lbl0_n_303, B2 => position_1(4), ZN => lbl0_n_335);
  lbl0_g14647 : ND2D1BWP7T port map(A1 => lbl0_n_322, A2 => lbl0_read_data_reg(0), ZN => lbl0_n_334);
  lbl0_g14648 : ND2D1BWP7T port map(A1 => lbl0_n_322, A2 => lbl0_read_data_reg(1), ZN => lbl0_n_333);
  lbl0_g14649 : OAI21D0BWP7T port map(A1 => lbl0_n_280, A2 => lbl0_n_294, B => lbl0_n_220, ZN => lbl0_d_position_0(1));
  lbl0_g14650 : OAI21D0BWP7T port map(A1 => lbl0_n_279, A2 => lbl0_n_296, B => lbl0_n_220, ZN => lbl0_d_position_1(1));
  lbl0_g14651 : NR2XD0BWP7T port map(A1 => lbl0_n_312, A2 => position_1(7), ZN => lbl0_n_341);
  lbl0_g14652 : AOI211XD0BWP7T port map(A1 => lbl0_n_269, A2 => position_0(2), B => lbl0_n_291, C => lbl0_n_275, ZN => lbl0_n_340);
  lbl0_g14653 : AOI22D0BWP7T port map(A1 => lbl0_n_276, A2 => lbl0_n_145, B1 => lbl0_next_direction_1(0), B2 => position_1(6), ZN => lbl0_n_339);
  lbl0_g14654 : AOI211XD0BWP7T port map(A1 => lbl0_n_270, A2 => position_1(2), B => lbl0_n_288, C => lbl0_n_141, ZN => lbl0_n_338);
  lbl0_g14655 : OAI21D0BWP7T port map(A1 => lbl0_n_299, A2 => lbl0_n_144, B => lbl0_n_300, ZN => lbl0_n_336);
  lbl0_g14656 : AOI22D0BWP7T port map(A1 => lbl0_n_301, A2 => position_0(3), B1 => lbl0_n_303, B2 => position_1(3), ZN => lbl0_n_329);
  lbl0_g14657 : AOI22D0BWP7T port map(A1 => lbl0_n_301, A2 => position_0(2), B1 => lbl0_n_303, B2 => position_1(2), ZN => lbl0_n_328);
  lbl0_g14658 : AOI22D0BWP7T port map(A1 => lbl0_n_301, A2 => position_0(0), B1 => lbl0_n_303, B2 => position_1(0), ZN => lbl0_n_327);
  lbl0_g14659 : AOI22D0BWP7T port map(A1 => lbl0_n_301, A2 => position_0(1), B1 => lbl0_n_303, B2 => position_1(1), ZN => lbl0_n_326);
  lbl0_g14660 : MOAI22D0BWP7T port map(A1 => lbl0_n_310, A2 => lbl0_next_layer_0, B1 => lbl0_n_142, B2 => lbl0_next_layer_0, ZN => lbl0_n_325);
  lbl0_g14661 : MOAI22D0BWP7T port map(A1 => lbl0_n_297, A2 => position_0(8), B1 => lbl0_n_297, B2 => position_0(8), ZN => lbl0_n_324);
  lbl0_g14662 : MOAI22D0BWP7T port map(A1 => lbl0_n_310, A2 => lbl0_next_layer_1, B1 => lbl0_n_142, B2 => lbl0_next_layer_1, ZN => lbl0_n_323);
  lbl0_g14663 : MAOI22D0BWP7T port map(A1 => lbl0_n_238, A2 => lbl0_n_167, B1 => lbl0_n_238, B2 => lbl0_n_167, ZN => lbl0_n_332);
  lbl0_g14664 : MAOI22D0BWP7T port map(A1 => lbl0_n_308, A2 => position_0(3), B1 => lbl0_n_308, B2 => position_0(3), ZN => lbl0_n_331);
  lbl0_g14665 : MAOI22D0BWP7T port map(A1 => lbl0_n_309, A2 => position_1(3), B1 => lbl0_n_309, B2 => position_1(3), ZN => lbl0_n_330);
  lbl0_g14666 : INVD1BWP7T port map(I => lbl0_n_320, ZN => lbl0_n_321);
  lbl0_g14667 : INVD1BWP7T port map(I => lbl0_n_319, ZN => lbl0_n_318);
  lbl0_g14668 : INVD0BWP7T port map(I => lbl0_n_317, ZN => lbl0_n_316);
  lbl0_g14669 : INR2D1BWP7T port map(A1 => read_memory_in(0), B1 => lbl0_n_298, ZN => lbl0_d_read_data_reg(0));
  lbl0_g14670 : INR2D1BWP7T port map(A1 => read_memory_in(1), B1 => lbl0_n_298, ZN => lbl0_d_read_data_reg(1));
  lbl0_g14671 : INR2D1BWP7T port map(A1 => read_memory_in(2), B1 => lbl0_n_298, ZN => lbl0_d_read_data_reg(2));
  lbl0_g14672 : INR2D1BWP7T port map(A1 => read_memory_in(7), B1 => lbl0_n_298, ZN => lbl0_d_read_data_reg(7));
  lbl0_g14673 : INR2D1BWP7T port map(A1 => read_memory_in(6), B1 => lbl0_n_298, ZN => lbl0_d_read_data_reg(6));
  lbl0_g14674 : INR2D1BWP7T port map(A1 => read_memory_in(5), B1 => lbl0_n_298, ZN => lbl0_d_read_data_reg(5));
  lbl0_g14675 : INR2D1BWP7T port map(A1 => read_memory_in(4), B1 => lbl0_n_298, ZN => lbl0_d_read_data_reg(4));
  lbl0_g14676 : INR2D1BWP7T port map(A1 => read_memory_in(3), B1 => lbl0_n_298, ZN => lbl0_d_read_data_reg(3));
  lbl0_g14677 : INR2D1BWP7T port map(A1 => lbl0_n_297, B1 => position_0(7), ZN => lbl0_n_315);
  lbl0_g14678 : ND2D1BWP7T port map(A1 => lbl0_n_306, A2 => lbl0_n_143, ZN => lbl0_n_322);
  lbl0_g14679 : ND2D1BWP7T port map(A1 => lbl0_n_304, A2 => lbl0_n_307, ZN => lbl0_n_320);
  lbl0_g14680 : NR2D1BWP7T port map(A1 => lbl0_n_302, A2 => lbl0_next_direction_1(0), ZN => lbl0_n_319);
  lbl0_g14681 : NR2D1BWP7T port map(A1 => lbl0_n_299, A2 => lbl0_next_direction_0(0), ZN => lbl0_n_317);
  lbl0_g14682 : MOAI22D0BWP7T port map(A1 => lbl0_n_278, A2 => position_0(10), B1 => lbl0_n_271, B2 => position_0(10), ZN => lbl0_n_472);
  lbl0_g14683 : MOAI22D0BWP7T port map(A1 => lbl0_n_273, A2 => position_1(10), B1 => lbl0_n_268, B2 => position_1(10), ZN => lbl0_n_471);
  lbl0_g14684 : OAI21D0BWP7T port map(A1 => lbl0_n_277, A2 => position_0(10), B => lbl0_n_290, ZN => lbl0_n_474);
  lbl0_g14685 : OAI21D0BWP7T port map(A1 => lbl0_n_272, A2 => position_1(10), B => lbl0_n_289, ZN => lbl0_n_473);
  lbl0_g14686 : MOAI22D0BWP7T port map(A1 => lbl0_n_279, A2 => lbl0_n_204, B1 => lbl0_n_505, B2 => start_position_1(5), ZN => lbl0_d_position_1(5));
  lbl0_g14687 : IOA21D1BWP7T port map(A1 => lbl0_n_281, A2 => FE_PHN59_lbl0_next_layer_0, B => lbl0_n_168, ZN => lbl0_d_layer_0);
  lbl0_g14688 : OAI21D0BWP7T port map(A1 => lbl0_n_279, A2 => FE_PHN61_lbl0_n_148, B => lbl0_n_168, ZN => lbl0_d_layer_1);
  lbl0_g14689 : OAI21D0BWP7T port map(A1 => lbl0_n_279, A2 => lbl0_n_200, B => lbl0_n_168, ZN => lbl0_d_position_1(0));
  lbl0_g14691 : MUX2ND0BWP7T port map(I0 => lbl0_n_141, I1 => lbl0_n_266, S => position_1(3), ZN => lbl0_n_314);
  lbl0_g14692 : MAOI22D0BWP7T port map(A1 => lbl0_n_286, A2 => lbl0_n_181, B1 => lbl0_n_286, B2 => lbl0_n_181, ZN => lbl0_n_313);
  lbl0_g14693 : IAO21D0BWP7T port map(A1 => lbl0_n_167, A2 => position_1(7), B => lbl0_n_238, ZN => lbl0_n_312);
  lbl0_g14694 : AOI22D0BWP7T port map(A1 => lbl0_n_287, A2 => lbl0_n_144, B1 => lbl0_next_direction_0(0), B2 => position_0(6), ZN => lbl0_n_311);
  lbl0_g14695 : INVD1BWP7T port map(I => lbl0_n_305, ZN => lbl0_n_304);
  lbl0_g14696 : INVD1BWP7T port map(I => lbl0_n_300, ZN => lbl0_n_301);
  lbl0_g14697 : NR2D1BWP7T port map(A1 => lbl0_n_280, A2 => lbl0_n_202, ZN => lbl0_n_413);
  lbl0_g14698 : OAI31D0BWP7T port map(A1 => read_memory_in(0), A2 => read_memory_in(1), A3 => lbl0_n_165, B => lbl0_n_283, ZN => lbl0_n_310);
  lbl0_g14699 : NR2XD0BWP7T port map(A1 => lbl0_n_141, A2 => lbl0_n_266, ZN => lbl0_n_309);
  lbl0_g14701 : NR2XD0BWP7T port map(A1 => lbl0_n_275, A2 => lbl0_n_265, ZN => lbl0_n_308);
  lbl0_g14702 : IND2D1BWP7T port map(A1 => position_0(10), B1 => lbl0_n_284, ZN => lbl0_n_307);
  lbl0_g14703 : ND2D1BWP7T port map(A1 => lbl0_n_284, A2 => position_0(10), ZN => lbl0_n_306);
  lbl0_g14705 : NR2XD0BWP7T port map(A1 => lbl0_n_285, A2 => position_1(10), ZN => lbl0_n_305);
  lbl0_g14706 : OA21D0BWP7T port map(A1 => lbl0_n_213, A2 => lbl0_n_225, B => lbl0_n_282, Z => lbl0_n_303);
  lbl0_g14707 : ND2D1BWP7T port map(A1 => lbl0_n_282, A2 => lbl0_n_227, ZN => lbl0_n_302);
  lbl0_g14708 : ND2D1BWP7T port map(A1 => lbl0_n_260, A2 => lbl0_n_282, ZN => lbl0_n_300);
  lbl0_g14709 : ND2D1BWP7T port map(A1 => lbl0_n_282, A2 => lbl0_n_241, ZN => lbl0_n_299);
  lbl0_g14710 : ND2D1BWP7T port map(A1 => lbl0_n_283, A2 => lbl0_n_430, ZN => lbl0_n_298);
  lbl0_g14711 : INVD1BWP7T port map(I => lbl0_n_295, ZN => lbl0_n_296);
  lbl0_g14712 : INVD1BWP7T port map(I => lbl0_n_293, ZN => lbl0_n_294);
  lbl0_g14713 : IOA21D1BWP7T port map(A1 => lbl0_n_504, A2 => FE_PHN58_lbl0_next_direction_0_1, B => lbl0_n_168, ZN => lbl0_d_direction_0(1));
  lbl0_g14714 : NR4D0BWP7T port map(A1 => lbl0_n_244, A2 => lbl0_n_508, A3 => lbl0_n_513, A4 => lbl0_n_417, ZN => lbl0_n_292);
  lbl0_g14715 : OAI31D0BWP7T port map(A1 => position_0(2), A2 => lbl0_n_183, A3 => lbl0_n_190, B => lbl0_n_139, ZN => lbl0_n_291);
  lbl0_g14716 : OAI21D0BWP7T port map(A1 => lbl0_n_232, A2 => lbl0_n_257, B => position_0(10), ZN => lbl0_n_290);
  lbl0_g14717 : OAI21D0BWP7T port map(A1 => lbl0_n_233, A2 => lbl0_n_250, B => position_1(10), ZN => lbl0_n_289);
  lbl0_g14718 : IOA21D1BWP7T port map(A1 => lbl0_n_504, A2 => lbl0_next_direction_1(0), B => lbl0_n_216, ZN => lbl0_d_direction_1(0));
  lbl0_g14719 : OAI31D0BWP7T port map(A1 => position_1(2), A2 => lbl0_n_169, A3 => lbl0_n_176, B => lbl0_n_140, ZN => lbl0_n_288);
  lbl0_g14720 : NR2D1BWP7T port map(A1 => lbl0_n_280, A2 => lbl0_n_205, ZN => lbl0_n_411);
  lbl0_g14721 : IOA21D1BWP7T port map(A1 => lbl0_n_504, A2 => lbl0_next_direction_0(0), B => lbl0_n_216, ZN => lbl0_d_direction_0(0));
  lbl0_g14722 : AOI21D1BWP7T port map(A1 => lbl0_n_504, A2 => lbl0_n_210, B => lbl0_n_236, ZN => lbl0_e_position_1);
  lbl0_g14723 : AOI21D1BWP7T port map(A1 => lbl0_n_504, A2 => lbl0_n_226, B => lbl0_n_236, ZN => lbl0_e_position_0);
  lbl0_g14724 : OAI221D1BWP7T port map(A1 => lbl0_n_192, A2 => lbl0_n_157, B1 => lbl0_mem_com_state(2), B2 => lbl0_n_177, C => lbl0_n_194, ZN => lbl0_n_427);
  lbl0_g14725 : OAI21D0BWP7T port map(A1 => lbl0_n_182, A2 => position_0(7), B => lbl0_n_286, ZN => lbl0_n_297);
  lbl0_g14726 : OAI21D0BWP7T port map(A1 => lbl0_n_134, A2 => lbl0_n_169, B => lbl0_n_274, ZN => lbl0_n_295);
  lbl0_g14727 : OAI21D0BWP7T port map(A1 => lbl0_n_136, A2 => lbl0_n_183, B => lbl0_n_267, ZN => lbl0_n_293);
  lbl0_g14730 : INVD1BWP7T port map(I => lbl0_n_281, ZN => lbl0_n_280);
  lbl0_g14731 : FA1D0BWP7T port map(A => position_0(5), B => position_0(6), CI => lbl0_n_182, CO => lbl0_n_286, S => lbl0_n_287);
  lbl0_g14732 : AN2D0BWP7T port map(A1 => lbl0_n_425, A2 => direction_in(0), Z => lbl0_d_next_direction_0(0));
  lbl0_g14733 : AOI221D0BWP7T port map(A1 => borders(0), A2 => lbl0_n_182, B1 => borders(1), B2 => lbl0_n_172, C => lbl0_n_255, ZN => lbl0_n_278);
  lbl0_g14734 : INR2D1BWP7T port map(A1 => lbl0_n_509, B1 => FE_PHN30_lbl0_booster_sync, ZN => lbl0_d_booster_sync);
  lbl0_g14735 : AN2D0BWP7T port map(A1 => lbl0_n_504, A2 => FE_PHN39_lbl0_next_direction_1_1, Z => lbl0_d_direction_1(1));
  lbl0_g14736 : AOI221D0BWP7T port map(A1 => lbl0_n_182, A2 => ramps(0), B1 => ramps(1), B2 => lbl0_n_172, C => lbl0_n_252, ZN => lbl0_n_277);
  lbl0_g14737 : OR2D1BWP7T port map(A1 => lbl0_n_509, A2 => lbl0_n_505, Z => lbl0_n_432);
  lbl0_g14738 : AN2D0BWP7T port map(A1 => lbl0_n_425, A2 => direction_in(1), Z => lbl0_d_next_direction_0(1));
  lbl0_g14739 : AN2D0BWP7T port map(A1 => lbl0_n_424, A2 => direction_in(2), Z => lbl0_d_next_direction_1(0));
  lbl0_g14740 : AN2D0BWP7T port map(A1 => lbl0_n_424, A2 => direction_in(3), Z => lbl0_d_next_direction_1(1));
  lbl0_g14741 : ND2D1BWP7T port map(A1 => lbl0_n_423, A2 => lbl0_n_225, ZN => lbl0_n_285);
  lbl0_g14742 : INR2XD0BWP7T port map(A1 => lbl0_n_423, B1 => lbl0_n_246, ZN => lbl0_n_284);
  lbl0_g14743 : NR3D0BWP7T port map(A1 => lbl0_n_198, A2 => lbl0_n_152, A3 => lbl0_mem_com_state(3), ZN => lbl0_n_283);
  lbl0_g14744 : AOI211XD0BWP7T port map(A1 => lbl0_n_174, A2 => lbl0_n_157, B => lbl0_n_214, C => lbl0_mem_com_state(3), ZN => lbl0_n_282);
  lbl0_g14745 : INR2XD0BWP7T port map(A1 => lbl0_n_504, B1 => lbl0_n_226, ZN => lbl0_n_281);
  lbl0_g14746 : IND2D1BWP7T port map(A1 => lbl0_n_210, B1 => lbl0_n_504, ZN => lbl0_n_279);
  lbl0_g14747 : AOI22D0BWP7T port map(A1 => lbl0_n_134, A2 => lbl0_n_185, B1 => lbl0_n_145, B2 => position_1(1), ZN => lbl0_n_274);
  lbl0_g14748 : AOI221D0BWP7T port map(A1 => borders(0), A2 => lbl0_n_167, B1 => borders(1), B2 => lbl0_n_185, C => lbl0_n_253, ZN => lbl0_n_273);
  lbl0_g14749 : AOI221D0BWP7T port map(A1 => lbl0_n_167, A2 => ramps(0), B1 => ramps(1), B2 => lbl0_n_185, C => lbl0_n_251, ZN => lbl0_n_272);
  lbl0_g14750 : ND2D1BWP7T port map(A1 => lbl0_n_235, A2 => lbl0_n_256, ZN => lbl0_n_271);
  lbl0_g14751 : AO21D0BWP7T port map(A1 => lbl0_n_174, A2 => lbl0_mem_com_state(1), B => lbl0_n_237, Z => write_enable);
  lbl0_g14752 : OAI21D0BWP7T port map(A1 => lbl0_n_186, A2 => lbl0_n_180, B => lbl0_next_direction_1(0), ZN => lbl0_n_270);
  lbl0_g14753 : OA21D0BWP7T port map(A1 => lbl0_n_138, A2 => FE_PHN30_lbl0_booster_sync, B => lbl0_n_509, Z => lbl0_d_booster_0);
  lbl0_g14754 : OA21D0BWP7T port map(A1 => lbl0_n_242, A2 => FE_PHN30_lbl0_booster_sync, B => lbl0_n_509, Z => lbl0_d_booster_1);
  lbl0_g14755 : OAI21D0BWP7T port map(A1 => lbl0_n_171, A2 => lbl0_n_195, B => lbl0_next_direction_0(0), ZN => lbl0_n_269);
  lbl0_g14756 : OAI211D1BWP7T port map(A1 => lbl0_state(1), A2 => lbl0_n_156, B => lbl0_n_247, C => lbl0_n_410, ZN => game_state(0));
  lbl0_g14757 : IIND4D0BWP7T port map(A1 => lbl0_n_436, A2 => lbl0_n_437, B1 => lbl0_n_410, B2 => lbl0_n_173, ZN => game_state(1));
  lbl0_g14758 : ND2D1BWP7T port map(A1 => lbl0_n_231, A2 => lbl0_n_254, ZN => lbl0_n_268);
  lbl0_g14759 : AOI22D0BWP7T port map(A1 => lbl0_n_136, A2 => lbl0_n_172, B1 => lbl0_n_144, B2 => position_0(1), ZN => lbl0_n_267);
  lbl0_g14760 : MOAI22D0BWP7T port map(A1 => lbl0_n_239, A2 => position_1(6), B1 => lbl0_n_239, B2 => position_1(6), ZN => lbl0_n_276);
  lbl0_g14761 : AN3D1BWP7T port map(A1 => lbl0_n_172, A2 => lbl0_n_195, A3 => lbl0_n_150, Z => lbl0_n_275);
  lbl0_g14763 : AN2D0BWP7T port map(A1 => lbl0_n_512, A2 => direction_in(2), Z => lbl0_d_speed_select(0));
  lbl0_g14764 : AN2D0BWP7T port map(A1 => lbl0_n_512, A2 => direction_in(3), Z => lbl0_d_speed_select(1));
  lbl0_g14765 : IND2D0BWP7T port map(A1 => lbl0_n_428, B1 => lbl0_n_511, ZN => lbl0_n_264);
  lbl0_g14766 : NR2XD0BWP7T port map(A1 => lbl0_n_177, A2 => lbl0_n_152, ZN => clear_memory);
  lbl0_g14767 : IND2D0BWP7T port map(A1 => lbl0_n_429, B1 => lbl0_n_511, ZN => lbl0_n_263);
  lbl0_g14768 : OR2D1BWP7T port map(A1 => lbl0_n_237, A2 => lbl0_mem_com_n_175, Z => go_to);
  lbl0_g14771 : NR2D1BWP7T port map(A1 => lbl0_n_230, A2 => lbl0_n_176, ZN => lbl0_n_266);
  lbl0_g14772 : NR2D1BWP7T port map(A1 => lbl0_n_228, A2 => lbl0_n_190, ZN => lbl0_n_265);
  lbl0_g14773 : INR2XD0BWP7T port map(A1 => lbl0_n_244, B1 => lbl0_n_242, ZN => lbl0_n_424);
  lbl0_g14774 : OR2D1BWP7T port map(A1 => lbl0_n_418, A2 => lbl0_n_237, Z => lbl0_n_423);
  lbl0_g14775 : OR2D1BWP7T port map(A1 => lbl0_n_513, A2 => lbl0_n_511, Z => lbl0_n_422);
  lbl0_g14776 : INR2XD0BWP7T port map(A1 => lbl0_n_244, B1 => lbl0_n_138, ZN => lbl0_n_425);
  lbl0_g14777 : AN2D1BWP7T port map(A1 => lbl0_n_426, A2 => lbl0_state(1), Z => lbl0_n_509);
  lbl0_g14778 : NR2D1BWP7T port map(A1 => lbl0_n_236, A2 => lbl0_state(3), ZN => lbl0_n_504);
  lbl0_g14779 : AN2D0BWP7T port map(A1 => lbl0_n_512, A2 => direction_in(1), Z => lbl0_d_map_select(1));
  lbl0_g14780 : AN2D0BWP7T port map(A1 => lbl0_n_512, A2 => direction_in(0), Z => lbl0_d_map_select(0));
  lbl0_g14781 : AN2D0BWP7T port map(A1 => lbl0_n_417, A2 => lbl0_n_156, Z => lbl0_n_510);
  lbl0_g14782 : ND2D1BWP7T port map(A1 => lbl0_n_247, A2 => lbl0_n_187, ZN => game_state(2));
  lbl0_g14783 : IOA21D1BWP7T port map(A1 => lbl0_n_430, A2 => lbl0_n_8, B => lbl0_n_246, ZN => lbl0_n_260);
  lbl0_g14784 : MOAI22D0BWP7T port map(A1 => lbl0_n_200, A2 => position_0(0), B1 => lbl0_n_200, B2 => position_0(0), ZN => lbl0_n_259);
  lbl0_g14785 : XNR2D1BWP7T port map(A1 => lbl0_n_205, A2 => lbl0_n_200, ZN => lbl0_n_258);
  lbl0_g14786 : OAI22D0BWP7T port map(A1 => lbl0_n_222, A2 => ramps(6), B1 => ramps(7), B2 => lbl0_n_183, ZN => lbl0_n_257);
  lbl0_g14787 : AOI22D0BWP7T port map(A1 => borders(6), A2 => lbl0_n_223, B1 => borders(7), B2 => lbl0_n_184, ZN => lbl0_n_256);
  lbl0_g14788 : AO22D0BWP7T port map(A1 => borders(2), A2 => lbl0_n_223, B1 => lbl0_n_184, B2 => borders(3), Z => lbl0_n_255);
  lbl0_g14789 : AOI22D0BWP7T port map(A1 => borders(6), A2 => lbl0_n_218, B1 => borders(7), B2 => lbl0_n_170, ZN => lbl0_n_254);
  lbl0_g14790 : AO22D0BWP7T port map(A1 => borders(2), A2 => lbl0_n_218, B1 => lbl0_n_170, B2 => borders(3), Z => lbl0_n_253);
  lbl0_g14791 : AO22D0BWP7T port map(A1 => lbl0_n_223, A2 => ramps(2), B1 => lbl0_n_184, B2 => ramps(3), Z => lbl0_n_252);
  lbl0_g14792 : AO22D0BWP7T port map(A1 => lbl0_n_218, A2 => ramps(2), B1 => lbl0_n_170, B2 => ramps(3), Z => lbl0_n_251);
  lbl0_g14793 : OAI22D0BWP7T port map(A1 => lbl0_n_217, A2 => ramps(6), B1 => ramps(7), B2 => lbl0_n_169, ZN => lbl0_n_250);
  lbl0_g14794 : OAI222D0BWP7T port map(A1 => lbl0_n_162, A2 => lbl0_next_direction_1(1), B1 => direction_1(0), B2 => lbl0_next_direction_1(0), C1 => direction_1(1), C2 => lbl0_n_149, ZN => lbl0_n_262);
  lbl0_g14795 : OAI222D0BWP7T port map(A1 => lbl0_n_161, A2 => lbl0_next_direction_0(1), B1 => direction_0(0), B2 => lbl0_next_direction_0(0), C1 => direction_0(1), C2 => lbl0_n_151, ZN => lbl0_n_261);
  lbl0_g14797 : INVD0BWP7T port map(I => lbl0_n_207, ZN => lbl0_n_249);
  lbl0_g14798 : NR2D1BWP7T port map(A1 => lbl0_n_229, A2 => lbl0_mem_com_state(1), ZN => lbl0_mem_com_n_166);
  lbl0_g14799 : AN2D1BWP7T port map(A1 => lbl0_n_224, A2 => lbl0_state(4), Z => lbl0_n_507);
  lbl0_g14800 : ND2D1BWP7T port map(A1 => lbl0_n_221, A2 => FE_PHN42_lbl0_border_1, ZN => lbl0_n_248);
  lbl0_g14801 : CKND2D1BWP7T port map(A1 => lbl0_n_212, A2 => lbl0_n_211, ZN => lbl0_n_429);
  lbl0_g14802 : CKND2D1BWP7T port map(A1 => lbl0_n_209, A2 => lbl0_n_206, ZN => lbl0_n_428);
  lbl0_g14803 : INR2XD0BWP7T port map(A1 => lbl0_n_197, B1 => lbl0_state(3), ZN => lbl0_n_247);
  lbl0_g14804 : NR2D1BWP7T port map(A1 => lbl0_n_219, A2 => lbl0_n_188, ZN => lbl0_n_508);
  lbl0_g14806 : ND2D1BWP7T port map(A1 => lbl0_n_224, A2 => lbl0_state(3), ZN => lbl0_n_246);
  lbl0_g14807 : ND2D1BWP7T port map(A1 => lbl0_n_221, A2 => FE_PHN51_lbl0_border_0, ZN => lbl0_n_245);
  lbl0_g14808 : NR2XD0BWP7T port map(A1 => lbl0_n_229, A2 => lbl0_n_157, ZN => lbl0_n_418);
  lbl0_g14809 : NR2D0BWP7T port map(A1 => lbl0_n_219, A2 => lbl0_n_187, ZN => lbl0_n_513);
  lbl0_g14810 : INR2D1BWP7T port map(A1 => lbl0_n_224, B1 => lbl0_state(3), ZN => lbl0_n_417);
  lbl0_g14811 : NR2D1BWP7T port map(A1 => lbl0_n_219, A2 => lbl0_n_173, ZN => lbl0_n_244);
  lbl0_g14812 : NR2D1BWP7T port map(A1 => lbl0_n_219, A2 => lbl0_n_419, ZN => lbl0_n_511);
  lbl0_g14813 : INVD0BWP7T port map(I => lbl0_n_433, ZN => lbl0_n_236);
  lbl0_g14814 : AOI22D0BWP7T port map(A1 => borders(4), A2 => lbl0_n_182, B1 => borders(5), B2 => lbl0_n_172, ZN => lbl0_n_235);
  lbl0_g14815 : NR4D0BWP7T port map(A1 => read_memory_in(7), A2 => read_memory_in(6), A3 => read_memory_in(5), A4 => read_memory_in(4), ZN => lbl0_n_234);
  lbl0_g14816 : OAI22D0BWP7T port map(A1 => ramps(4), A2 => lbl0_n_166, B1 => ramps(5), B2 => lbl0_n_186, ZN => lbl0_n_233);
  lbl0_g14817 : OAI22D0BWP7T port map(A1 => ramps(4), A2 => lbl0_n_181, B1 => ramps(5), B2 => lbl0_n_171, ZN => lbl0_n_232);
  lbl0_g14818 : AOI22D0BWP7T port map(A1 => borders(4), A2 => lbl0_n_167, B1 => borders(5), B2 => lbl0_n_185, ZN => lbl0_n_231);
  lbl0_g14819 : MAOI22D0BWP7T port map(A1 => lbl0_n_178, A2 => lbl0_n_191, B1 => lbl0_n_178, B2 => lbl0_n_191, ZN => lbl0_n_243);
  lbl0_g14820 : INR2XD0BWP7T port map(A1 => lbl0_n_206, B1 => lbl0_n_209, ZN => lbl0_n_242);
  lbl0_g14821 : NR3D0BWP7T port map(A1 => lbl0_n_188, A2 => lbl0_n_147, A3 => lbl0_state(0), ZN => lbl0_n_241);
  lbl0_g14822 : MAOI22D0BWP7T port map(A1 => lbl0_n_179, A2 => lbl0_n_193, B1 => lbl0_n_179, B2 => lbl0_n_193, ZN => lbl0_n_240);
  lbl0_g14823 : MAOI22D0BWP7T port map(A1 => lbl0_n_166, A2 => position_1(5), B1 => lbl0_n_166, B2 => position_1(5), ZN => lbl0_n_239);
  lbl0_g14824 : MAOI222D1BWP7T port map(A => lbl0_n_167, B => position_1(6), C => position_1(5), ZN => lbl0_n_238);
  lbl0_g14825 : NR4D0BWP7T port map(A1 => lbl0_n_160, A2 => lbl0_mem_com_state(3), A3 => lbl0_mem_com_state(2), A4 => lbl0_mem_com_state(1), ZN => lbl0_n_237);
  lbl0_g14826 : NR3D0BWP7T port map(A1 => lbl0_n_189, A2 => lbl0_state(2), A3 => lbl0_state(0), ZN => lbl0_n_426);
  lbl0_g14827 : NR3D0BWP7T port map(A1 => lbl0_n_187, A2 => lbl0_n_156, A3 => lbl0_state(0), ZN => lbl0_n_433);
  lbl0_g14828 : NR3D1BWP7T port map(A1 => lbl0_n_189, A2 => lbl0_n_419, A3 => lbl0_state(0), ZN => lbl0_n_512);
  lbl0_g14831 : INVD0BWP7T port map(I => lbl0_n_223, ZN => lbl0_n_222);
  lbl0_g14832 : INVD0BWP7T port map(I => lbl0_n_218, ZN => lbl0_n_217);
  lbl0_g14833 : INVD1BWP7T port map(I => lbl0_n_215, ZN => lbl0_n_216);
  lbl0_g14834 : NR2D1BWP7T port map(A1 => lbl0_n_174, A2 => lbl0_n_157, ZN => lbl0_n_214);
  lbl0_g14836 : NR2D1BWP7T port map(A1 => lbl0_n_187, A2 => lbl0_n_175, ZN => lbl0_n_213);
  lbl0_g14837 : NR2D1BWP7T port map(A1 => lbl0_n_173, A2 => lbl0_n_410, ZN => lbl0_n_506);
  lbl0_g14838 : ND2D1BWP7T port map(A1 => lbl0_n_170, A2 => position_1(2), ZN => lbl0_n_230);
  lbl0_g14839 : IND2D1BWP7T port map(A1 => lbl0_mem_com_state(3), B1 => lbl0_n_174, ZN => lbl0_n_229);
  lbl0_g14840 : NR2XD0BWP7T port map(A1 => lbl0_n_192, A2 => lbl0_mem_com_state(1), ZN => lbl0_mem_com_n_175);
  lbl0_g14841 : ND2D1BWP7T port map(A1 => lbl0_n_184, A2 => position_0(2), ZN => lbl0_n_228);
  lbl0_g14842 : NR2XD0BWP7T port map(A1 => lbl0_n_188, A2 => lbl0_n_175, ZN => lbl0_n_227);
  lbl0_g14843 : OAI21D0BWP7T port map(A1 => lbl0_n_154, A2 => player_state_0(1), B => lbl0_booster_0, ZN => lbl0_n_226);
  lbl0_g14844 : NR2XD0BWP7T port map(A1 => lbl0_n_173, A2 => lbl0_n_175, ZN => lbl0_n_225);
  lbl0_g14845 : INR2XD0BWP7T port map(A1 => lbl0_n_437, B1 => lbl0_n_187, ZN => lbl0_n_430);
  lbl0_g14846 : NR2D1BWP7T port map(A1 => lbl0_n_173, A2 => lbl0_state(0), ZN => lbl0_n_224);
  lbl0_g14847 : NR2D1BWP7T port map(A1 => lbl0_n_182, A2 => lbl0_next_direction_0(0), ZN => lbl0_n_223);
  lbl0_g14848 : NR2XD0BWP7T port map(A1 => lbl0_n_187, A2 => lbl0_n_410, ZN => lbl0_n_221);
  lbl0_g14849 : ND2D1BWP7T port map(A1 => start_position_0(2), A2 => lbl0_n_505, ZN => lbl0_n_220);
  lbl0_g14850 : OR2D1BWP7T port map(A1 => lbl0_n_189, A2 => lbl0_n_8, Z => lbl0_n_219);
  lbl0_g14851 : NR2D1BWP7T port map(A1 => lbl0_n_167, A2 => lbl0_next_direction_1(0), ZN => lbl0_n_218);
  lbl0_g14852 : NR2D1BWP7T port map(A1 => start_position_0(2), A2 => lbl0_n_168, ZN => lbl0_n_215);
  lbl0_g14854 : INVD0BWP7T port map(I => lbl0_n_204, ZN => lbl0_n_203);
  lbl0_g14855 : INVD0BWP7T port map(I => lbl0_n_202, ZN => lbl0_n_201);
  lbl0_g14856 : MOAI22D0BWP7T port map(A1 => lbl0_next_layer_0, A2 => lbl0_next_layer_1, B1 => lbl0_next_layer_1, B2 => lbl0_next_layer_0, ZN => lbl0_n_199);
  lbl0_g14857 : OAI21D0BWP7T port map(A1 => lbl0_mem_com_state(0), A2 => lbl0_mem_com_state(1), B => lbl0_n_177, ZN => lbl0_n_198);
  lbl0_g14858 : OAI21D0BWP7T port map(A1 => lbl0_state(0), A2 => lbl0_state(1), B => lbl0_state(2), ZN => lbl0_n_197);
  lbl0_g14860 : MAOI22D0BWP7T port map(A1 => lbl0_n_148, A2 => position_0(10), B1 => lbl0_n_148, B2 => position_0(10), ZN => lbl0_n_196);
  lbl0_g14861 : MOAI22D0BWP7T port map(A1 => direction_0(1), A2 => direction_in(1), B1 => direction_0(1), B2 => direction_in(1), ZN => lbl0_n_212);
  lbl0_g14863 : NR3D0BWP7T port map(A1 => lbl0_n_156, A2 => lbl0_state(3), A3 => lbl0_state(2), ZN => lbl0_n_436);
  lbl0_g14864 : MOAI22D0BWP7T port map(A1 => direction_0(0), A2 => direction_in(0), B1 => direction_0(0), B2 => direction_in(0), ZN => lbl0_n_211);
  lbl0_g14865 : OAI21D0BWP7T port map(A1 => lbl0_n_153, A2 => player_state_1(1), B => lbl0_booster_1, ZN => lbl0_n_210);
  lbl0_g14866 : MOAI22D0BWP7T port map(A1 => direction_1(1), A2 => direction_in(3), B1 => direction_1(1), B2 => direction_in(3), ZN => lbl0_n_209);
  lbl0_g14867 : MAOI22D0BWP7T port map(A1 => lbl0_n_144, A2 => direction_0(0), B1 => lbl0_n_144, B2 => direction_0(0), ZN => lbl0_n_208);
  lbl0_g14868 : MOAI22D0BWP7T port map(A1 => lbl0_n_145, A2 => direction_1(0), B1 => lbl0_n_145, B2 => direction_1(0), ZN => lbl0_n_207);
  lbl0_g14869 : MOAI22D0BWP7T port map(A1 => direction_1(0), A2 => direction_in(2), B1 => direction_1(0), B2 => direction_in(2), ZN => lbl0_n_206);
  lbl0_g14871 : MAOI22D0BWP7T port map(A1 => lbl0_n_144, A2 => position_0(0), B1 => lbl0_n_144, B2 => position_0(0), ZN => lbl0_n_205);
  lbl0_g14872 : MAOI22D0BWP7T port map(A1 => lbl0_next_direction_1(0), A2 => position_1(5), B1 => lbl0_next_direction_1(0), B2 => position_1(5), ZN => lbl0_n_204);
  lbl0_g14873 : MAOI22D0BWP7T port map(A1 => lbl0_next_direction_0(0), A2 => position_0(5), B1 => lbl0_next_direction_0(0), B2 => position_0(5), ZN => lbl0_n_202);
  lbl0_g14874 : MAOI22D0BWP7T port map(A1 => lbl0_n_145, A2 => position_1(0), B1 => lbl0_n_145, B2 => position_1(0), ZN => lbl0_n_200);
  lbl0_g14876 : INVD1BWP7T port map(I => lbl0_n_186, ZN => lbl0_n_185);
  lbl0_g14877 : INVD0BWP7T port map(I => lbl0_n_184, ZN => lbl0_n_183);
  lbl0_g14878 : INVD1BWP7T port map(I => lbl0_n_182, ZN => lbl0_n_181);
  lbl0_g14879 : CKND2D0BWP7T port map(A1 => lbl0_state(4), A2 => lbl0_state(2), ZN => lbl0_n_1952_BAR);
  lbl0_g14880 : NR2D1BWP7T port map(A1 => position_0(0), A2 => position_0(1), ZN => lbl0_n_195);
  lbl0_g14881 : ND2D1BWP7T port map(A1 => lbl0_mem_com_state(3), A2 => lbl0_mem_com_state(0), ZN => lbl0_n_194);
  lbl0_g14882 : IND2D1BWP7T port map(A1 => direction_0(0), B1 => lbl0_next_direction_0(1), ZN => lbl0_n_193);
  lbl0_g14883 : ND2D1BWP7T port map(A1 => lbl0_n_160, A2 => lbl0_mem_com_state(2), ZN => lbl0_n_192);
  lbl0_g14884 : IND2D1BWP7T port map(A1 => direction_1(0), B1 => lbl0_next_direction_1(1), ZN => lbl0_n_191);
  lbl0_g14885 : CKND2D1BWP7T port map(A1 => position_0(1), A2 => position_0(0), ZN => lbl0_n_190);
  lbl0_g14886 : ND2D1BWP7T port map(A1 => lbl0_n_156, A2 => lbl0_n_147, ZN => lbl0_n_189);
  lbl0_g14887 : IND2D1BWP7T port map(A1 => lbl0_state(2), B1 => lbl0_state(1), ZN => lbl0_n_188);
  lbl0_g14888 : IND2D1BWP7T port map(A1 => lbl0_state(1), B1 => lbl0_state(2), ZN => lbl0_n_419);
  lbl0_g14889 : OR2D1BWP7T port map(A1 => lbl0_state(2), A2 => lbl0_state(1), Z => lbl0_n_187);
  lbl0_g14890 : ND2D1BWP7T port map(A1 => lbl0_next_direction_1(0), A2 => lbl0_n_149, ZN => lbl0_n_186);
  lbl0_g14891 : NR2XD0BWP7T port map(A1 => lbl0_n_144, A2 => lbl0_n_151, ZN => lbl0_n_184);
  lbl0_g14892 : NR2XD0BWP7T port map(A1 => lbl0_next_direction_0(0), A2 => lbl0_next_direction_0(1), ZN => lbl0_n_182);
  lbl0_g14893 : INVD0BWP7T port map(I => lbl0_n_172, ZN => lbl0_n_171);
  lbl0_g14894 : INVD0BWP7T port map(I => lbl0_n_170, ZN => lbl0_n_169);
  lbl0_g14895 : INVD1BWP7T port map(I => lbl0_n_168, ZN => lbl0_n_505);
  lbl0_g14896 : INVD0BWP7T port map(I => lbl0_n_167, ZN => lbl0_n_166);
  lbl0_g14897 : OR2D1BWP7T port map(A1 => read_memory_in(2), A2 => read_memory_in(3), Z => lbl0_n_165);
  lbl0_g14898 : NR2XD0BWP7T port map(A1 => position_1(0), A2 => position_1(1), ZN => lbl0_n_180);
  lbl0_g14899 : NR2XD0BWP7T port map(A1 => lbl0_next_direction_0(0), A2 => direction_0(1), ZN => lbl0_n_179);
  lbl0_g14900 : NR2D1BWP7T port map(A1 => lbl0_next_direction_1(0), A2 => direction_1(1), ZN => lbl0_n_178);
  lbl0_g14901 : ND2D1BWP7T port map(A1 => lbl0_mem_com_state(1), A2 => lbl0_mem_com_state(0), ZN => lbl0_n_177);
  lbl0_g14902 : CKND2D1BWP7T port map(A1 => position_1(1), A2 => position_1(0), ZN => lbl0_n_176);
  lbl0_g14903 : ND2D1BWP7T port map(A1 => lbl0_state(3), A2 => lbl0_state(0), ZN => lbl0_n_175);
  lbl0_g14904 : NR2D1BWP7T port map(A1 => lbl0_n_147, A2 => lbl0_state(4), ZN => lbl0_n_437);
  lbl0_g14905 : NR2XD0BWP7T port map(A1 => lbl0_mem_com_state(2), A2 => lbl0_mem_com_state(0), ZN => lbl0_n_174);
  lbl0_g14906 : ND2D1BWP7T port map(A1 => lbl0_state(4), A2 => lbl0_state(0), ZN => lbl0_n_410);
  lbl0_g14907 : ND2D1BWP7T port map(A1 => lbl0_state(2), A2 => lbl0_state(1), ZN => lbl0_n_173);
  lbl0_g14908 : NR2XD0BWP7T port map(A1 => lbl0_n_144, A2 => lbl0_next_direction_0(1), ZN => lbl0_n_172);
  lbl0_g14909 : NR2XD0BWP7T port map(A1 => lbl0_n_145, A2 => lbl0_n_149, ZN => lbl0_n_170);
  lbl0_g14910 : ND2D1BWP7T port map(A1 => lbl0_state(4), A2 => lbl0_state(3), ZN => lbl0_n_168);
  lbl0_g14911 : NR2XD0BWP7T port map(A1 => lbl0_next_direction_1(0), A2 => lbl0_next_direction_1(1), ZN => lbl0_n_167);
  lbl0_g14912 : INVD0BWP7T port map(I => lbl0_read_data_reg(7), ZN => lbl0_n_164);
  lbl0_g14913 : INVD0BWP7T port map(I => lbl0_read_data_reg(5), ZN => lbl0_n_163);
  lbl0_g14914 : INVD0BWP7T port map(I => direction_1(1), ZN => lbl0_n_162);
  lbl0_g14915 : INVD0BWP7T port map(I => direction_0(1), ZN => lbl0_n_161);
  lbl0_g14920 : INVD0BWP7T port map(I => position_0(8), ZN => lbl0_n_159);
  lbl0_g14921 : INVD1BWP7T port map(I => position_1(8), ZN => lbl0_n_158);
  lbl0_g14924 : INVD0BWP7T port map(I => lbl0_read_data_reg(4), ZN => lbl0_n_155);
  lbl0_g14925 : CKND1BWP7T port map(I => player_state_0(0), ZN => lbl0_n_154);
  lbl0_g14926 : CKND1BWP7T port map(I => player_state_1(0), ZN => lbl0_n_153);
  lbl0_g14928 : INVD0BWP7T port map(I => lbl0_next_direction_0(1), ZN => lbl0_n_151);
  lbl0_g14931 : INVD0BWP7T port map(I => position_0(2), ZN => lbl0_n_150);
  lbl0_g14932 : INVD1BWP7T port map(I => lbl0_next_direction_1(1), ZN => lbl0_n_149);
  lbl0_g14933 : INVD0BWP7T port map(I => lbl0_next_layer_1, ZN => lbl0_n_148);
  lbl0_g14938 : INVD1BWP7T port map(I => lbl0_next_direction_1(0), ZN => lbl0_n_145);
  lbl0_g14939 : INVD1BWP7T port map(I => lbl0_next_direction_0(0), ZN => lbl0_n_144);
  lbl0_g2 : IND2D1BWP7T port map(A1 => lbl0_n_285, B1 => position_1(10), ZN => lbl0_n_143);
  lbl0_g14940 : INR2D1BWP7T port map(A1 => lbl0_n_283, B1 => lbl0_n_234, ZN => lbl0_n_142);
  lbl0_g14941 : INR3D0BWP7T port map(A1 => lbl0_n_180, B1 => lbl0_n_186, B2 => position_1(2), ZN => lbl0_n_141);
  lbl0_g14942 : IND2D1BWP7T port map(A1 => lbl0_n_230, B1 => lbl0_n_176, ZN => lbl0_n_140);
  lbl0_g14943 : IND2D1BWP7T port map(A1 => lbl0_n_228, B1 => lbl0_n_190, ZN => lbl0_n_139);
  lbl0_g14944 : INR2D1BWP7T port map(A1 => lbl0_n_211, B1 => lbl0_n_212, ZN => lbl0_n_138);
  lbl0_g14945 : MUX2ND0BWP7T port map(I0 => lbl0_n_275, I1 => lbl0_n_265, S => position_0(3), ZN => lbl0_n_137);
  lbl0_g14946 : XNR2D1BWP7T port map(A1 => position_0(0), A2 => position_0(1), ZN => lbl0_n_136);
  lbl0_g14947 : XNR2D1BWP7T port map(A1 => lbl0_next_layer_0, A2 => position_1(10), ZN => lbl0_n_135);
  lbl0_g14948 : XNR2D1BWP7T port map(A1 => position_1(0), A2 => position_1(1), ZN => lbl0_n_134);
  lbl0_counter_busy_counter_state_reg_0 : DFQD1BWP7T port map(CP => CTS_11, D => lbl0_n_63, Q => FE_PHN56_lbl0_counter_busy_counter_state_0);
  lbl0_counter_busy_counter_state_reg_1 : DFQD1BWP7T port map(CP => CTS_11, D => lbl0_n_83, Q => FE_PHN62_lbl0_counter_busy_counter_state_1);
  lbl0_counter_unsigned_busy_count_reg_1 : DFQD1BWP7T port map(CP => CTS_11, D => FE_PHN70_lbl0_n_106, Q => FE_PHN49_lbl0_unsigned_busy_count_1);
  lbl0_counter_unsigned_busy_count_reg_2 : DFQD1BWP7T port map(CP => CTS_11, D => lbl0_n_109, Q => lbl0_unsigned_busy_count(2));
  lbl0_counter_unsigned_busy_count_reg_3 : DFQD1BWP7T port map(CP => CTS_11, D => lbl0_n_108, Q => FE_PHN54_lbl0_unsigned_busy_count_3);
  lbl0_counter_unsigned_busy_count_reg_4 : DFQD1BWP7T port map(CP => CTS_11, D => FE_PHN67_lbl0_n_107, Q => lbl0_unsigned_busy_count(4));
  lbl0_counter_unsigned_busy_count_reg_5 : DFQD1BWP7T port map(CP => CTS_11, D => FE_PHN65_lbl0_n_117, Q => lbl0_unsigned_busy_count(5));
  lbl0_counter_unsigned_busy_count_reg_6 : DFQD1BWP7T port map(CP => CTS_11, D => lbl0_n_119, Q => FE_PHN57_lbl0_unsigned_busy_count_6);
  lbl0_mem_com_state_reg_3 : DFQD1BWP7T port map(CP => CTS_12, D => FE_PHN77_lbl0_n_91, Q => lbl0_mem_com_state(3));
  lbl0_state_reg_2 : DFQD1BWP7T port map(CP => CTS_11, D => lbl0_n_120, Q => lbl0_state(2));
  lbl0_g10992 : ND4D0BWP7T port map(A1 => lbl0_n_130, A2 => lbl0_n_1, A3 => lbl0_n_0, A4 => lbl0_n_48, ZN => lbl0_n_133);
  lbl0_g10993 : IND4D0BWP7T port map(A1 => lbl0_n_96, B1 => lbl0_n_48, B2 => lbl0_n_67, B3 => lbl0_n_128, ZN => lbl0_n_132);
  lbl0_g10996 : ND4D0BWP7T port map(A1 => lbl0_n_125, A2 => lbl0_n_1, A3 => lbl0_n_34, A4 => lbl0_n_49, ZN => lbl0_n_131);
  lbl0_g10997 : NR3D0BWP7T port map(A1 => lbl0_n_126, A2 => lbl0_n_35, A3 => lbl0_n_95, ZN => lbl0_n_130);
  lbl0_g10998 : IND4D0BWP7T port map(A1 => lbl0_n_124, B1 => lbl0_n_73, B2 => lbl0_n_67, B3 => lbl0_n_0, ZN => lbl0_n_129);
  lbl0_g10999 : OA221D0BWP7T port map(A1 => lbl0_n_78, A2 => lbl0_n_55, B1 => FE_PHN46_lbl0_booster_1, B2 => lbl0_n_73, C => lbl0_n_127, Z => lbl0_n_128);
  lbl0_g11000 : AOI22D0BWP7T port map(A1 => lbl0_n_123, A2 => FE_DBTN4_rst, B1 => lbl0_n_47, B2 => lbl0_state(1), ZN => lbl0_n_127);
  lbl0_g11001 : OAI22D0BWP7T port map(A1 => lbl0_n_121, A2 => lbl0_state(1), B1 => lbl0_n_49, B2 => lbl0_n_17, ZN => lbl0_n_126);
  lbl0_g11003 : NR4D0BWP7T port map(A1 => lbl0_n_115, A2 => lbl0_n_43, A3 => lbl0_n_37, A4 => lbl0_n_104, ZN => lbl0_n_125);
  lbl0_g11004 : OAI222D0BWP7T port map(A1 => lbl0_n_55, A2 => lbl0_n_76, B1 => lbl0_n_65, B2 => lbl0_n_114, C1 => FE_OFN3_rst, C2 => lbl0_n_85, ZN => lbl0_n_124);
  lbl0_g11007 : IND3D1BWP7T port map(A1 => lbl0_n_509, B1 => lbl0_n_41, B2 => lbl0_n_113, ZN => lbl0_n_123);
  lbl0_g11008 : IND4D0BWP7T port map(A1 => lbl0_n_516, B1 => lbl0_n_39, B2 => lbl0_n_105, B3 => lbl0_n_92, ZN => lbl0_n_122);
  lbl0_g11009 : MAOI22D0BWP7T port map(A1 => lbl0_n_436, A2 => lbl0_n_25, B1 => lbl0_n_116, B2 => lbl0_n_65, ZN => lbl0_n_121);
  lbl0_g11011 : OR4D1BWP7T port map(A1 => lbl0_n_89, A2 => lbl0_n_96, A3 => lbl0_n_90, A4 => lbl0_n_79, Z => lbl0_n_120);
  lbl0_g11012 : OAI31D0BWP7T port map(A1 => lbl0_unsigned_busy_count(6), A2 => lbl0_n_86, A3 => lbl0_n_72, B => lbl0_n_118, ZN => FE_PHN66_lbl0_n_119);
  lbl0_g11013 : OAI21D0BWP7T port map(A1 => lbl0_n_97, A2 => lbl0_n_54, B => lbl0_unsigned_busy_count(6), ZN => lbl0_n_118);
  lbl0_g11019 : OAI31D0BWP7T port map(A1 => lbl0_unsigned_busy_count(5), A2 => lbl0_n_64, A3 => lbl0_n_72, B => lbl0_n_112, ZN => lbl0_n_117);
  lbl0_g11020 : IAO21D0BWP7T port map(A1 => lbl0_n_102, A2 => test_button, B => lbl0_n_87, ZN => lbl0_n_116);
  lbl0_g11021 : OAI211D1BWP7T port map(A1 => FE_OFN3_rst, A2 => lbl0_n_46, B => lbl0_n_111, C => lbl0_n_81, ZN => lbl0_n_115);
  lbl0_g11022 : AOI22D0BWP7T port map(A1 => lbl0_n_102, A2 => lbl0_n_29, B1 => lbl0_n_88, B2 => test_button, ZN => lbl0_n_114);
  lbl0_g11023 : AOI22D0BWP7T port map(A1 => lbl0_n_103, A2 => lbl0_n_510, B1 => lbl0_n_22, B2 => lbl0_n_14, ZN => lbl0_n_113);
  lbl0_g11025 : OAI21D0BWP7T port map(A1 => lbl0_n_84, A2 => lbl0_n_54, B => lbl0_unsigned_busy_count(5), ZN => lbl0_n_112);
  lbl0_g11026 : MAOI22D0BWP7T port map(A1 => lbl0_n_80, A2 => lbl0_state(1), B1 => lbl0_n_40, B2 => lbl0_n_10, ZN => lbl0_n_111);
  lbl0_g11027 : ND2D1BWP7T port map(A1 => lbl0_n_93, A2 => lbl0_n_39, ZN => FE_PHN75_lbl0_n_110);
  lbl0_g11030 : OAI31D0BWP7T port map(A1 => FE_PHN50_lbl0_unsigned_busy_count_2, A2 => lbl0_n_16, A3 => lbl0_n_72, B => lbl0_n_98, ZN => lbl0_n_109);
  lbl0_g11031 : OAI31D0BWP7T port map(A1 => FE_PHN80_lbl0_unsigned_busy_count_3, A2 => lbl0_n_38, A3 => lbl0_n_72, B => lbl0_n_100, ZN => lbl0_n_108);
  lbl0_g11032 : OAI31D0BWP7T port map(A1 => lbl0_unsigned_busy_count(4), A2 => lbl0_n_58, A3 => lbl0_n_72, B => lbl0_n_101, ZN => lbl0_n_107);
  lbl0_g11033 : OAI31D0BWP7T port map(A1 => lbl0_unsigned_busy_count(1), A2 => lbl0_n_7, A3 => lbl0_n_72, B => lbl0_n_99, ZN => lbl0_n_106);
  lbl0_g11034 : AOI22D0BWP7T port map(A1 => memory_ready, A2 => lbl0_n_82, B1 => lbl0_mem_com_n_175, B2 => lbl0_n_18, ZN => lbl0_n_105);
  lbl0_g11035 : AO33D0BWP7T port map(A1 => lbl0_n_427, A2 => lbl0_n_74, A3 => lbl0_n_17, B1 => lbl0_n_44, B2 => lbl0_n_437, B3 => lbl0_n_4, Z => lbl0_n_104);
  lbl0_g11037 : OAI21D0BWP7T port map(A1 => lbl0_n_68, A2 => lbl0_n_54, B => lbl0_unsigned_busy_count(4), ZN => lbl0_n_101);
  lbl0_g11038 : OAI21D0BWP7T port map(A1 => lbl0_n_61, A2 => lbl0_n_54, B => lbl0_unsigned_busy_count(3), ZN => lbl0_n_100);
  lbl0_g11039 : OAI21D0BWP7T port map(A1 => lbl0_n_70, A2 => lbl0_n_54, B => lbl0_unsigned_busy_count(1), ZN => lbl0_n_99);
  lbl0_g11040 : OAI21D0BWP7T port map(A1 => lbl0_n_71, A2 => lbl0_n_54, B => FE_PHN50_lbl0_unsigned_busy_count_2, ZN => lbl0_n_98);
  lbl0_g11041 : INR2D1BWP7T port map(A1 => lbl0_n_86, B1 => lbl0_n_53, ZN => lbl0_n_97);
  lbl0_g11042 : IND2D1BWP7T port map(A1 => lbl0_n_86, B1 => lbl0_unsigned_busy_count(6), ZN => lbl0_n_103);
  lbl0_g11043 : AOI221D0BWP7T port map(A1 => lbl0_n_51, A2 => lbl0_unsigned_busy_count(3), B1 => lbl0_n_52, B2 => FE_PHN50_lbl0_unsigned_busy_count_2, C => lbl0_unsigned_busy_count(4), ZN => lbl0_n_102);
  lbl0_g11045 : OAI32D1BWP7T port map(A1 => lbl0_n_10, A2 => lbl0_n_14, A3 => lbl0_n_21, B1 => lbl0_n_75, B2 => lbl0_n_55, ZN => lbl0_n_95);
  lbl0_g11046 : MOAI22D0BWP7T port map(A1 => lbl0_n_72, A2 => lbl0_unsigned_busy_count(0), B1 => lbl0_n_54, B2 => lbl0_unsigned_busy_count(0), ZN => lbl0_n_94);
  lbl0_g11047 : AOI32D1BWP7T port map(A1 => memory_ready, A2 => lbl0_n_57, A3 => FE_PHN36_lbl0_mem_com_state_0, B1 => lbl0_n_423, B2 => FE_DBTN4_rst, ZN => lbl0_n_93);
  lbl0_g11048 : AOI22D0BWP7T port map(A1 => lbl0_n_69, A2 => FE_PHN36_lbl0_mem_com_state_0, B1 => lbl0_mem_com_n_166, B2 => lbl0_n_50, ZN => lbl0_n_92);
  lbl0_g11049 : AO211D0BWP7T port map(A1 => clear_memory, A2 => lbl0_n_18, B => lbl0_n_516, C => lbl0_n_66, Z => lbl0_n_91);
  lbl0_g11050 : AO221D0BWP7T port map(A1 => lbl0_n_15, A2 => lbl0_n_427, B1 => lbl0_n_22, B2 => lbl0_n_515, C => lbl0_n_31, Z => lbl0_n_90);
  lbl0_g11051 : MOAI22D0BWP7T port map(A1 => lbl0_n_55, A2 => lbl0_n_77, B1 => lbl0_n_47, B2 => lbl0_n_4, ZN => lbl0_n_89);
  lbl0_g11052 : AO21D0BWP7T port map(A1 => lbl0_n_5, A2 => lbl0_n_74, B => lbl0_n_35, Z => lbl0_n_96);
  lbl0_g11053 : INVD0BWP7T port map(I => lbl0_n_87, ZN => lbl0_n_88);
  lbl0_g11054 : INR3D0BWP7T port map(A1 => lbl0_n_45, B1 => lbl0_n_504, B2 => lbl0_n_508, ZN => lbl0_n_85);
  lbl0_g11055 : INR2XD0BWP7T port map(A1 => lbl0_n_64, B1 => lbl0_n_53, ZN => lbl0_n_84);
  lbl0_g11056 : ND2D1BWP7T port map(A1 => lbl0_n_64, A2 => lbl0_n_29, ZN => lbl0_n_87);
  lbl0_g11057 : IND2D1BWP7T port map(A1 => lbl0_n_64, B1 => lbl0_unsigned_busy_count(5), ZN => lbl0_n_86);
  lbl0_g11060 : OAI22D0BWP7T port map(A1 => lbl0_n_36, A2 => lbl0_n_32, B1 => lbl0_n_53, B2 => lbl0_counter_busy_counter_state(0), ZN => lbl0_n_83);
  lbl0_g11061 : AO21D0BWP7T port map(A1 => lbl0_n_418, A2 => FE_DBTN4_rst, B => lbl0_n_66, Z => lbl0_n_82);
  lbl0_g11062 : IOA21D1BWP7T port map(A1 => lbl0_n_48, A2 => lbl0_n_517, B => lbl0_state(0), ZN => lbl0_n_81);
  lbl0_g11063 : AOI21D0BWP7T port map(A1 => lbl0_n_427, A2 => lbl0_booster_0, B => lbl0_n_65, ZN => lbl0_n_80);
  lbl0_g11064 : OAI22D0BWP7T port map(A1 => lbl0_n_60, A2 => lbl0_n_10, B1 => lbl0_n_34, B2 => FE_PHN46_lbl0_booster_1, ZN => lbl0_n_79);
  lbl0_g11066 : INVD0BWP7T port map(I => lbl0_n_77, ZN => lbl0_n_78);
  lbl0_g11067 : CKND1BWP7T port map(I => lbl0_n_75, ZN => lbl0_n_76);
  lbl0_g11068 : INVD0BWP7T port map(I => lbl0_n_74, ZN => lbl0_n_73);
  lbl0_g11069 : HA1D0BWP7T port map(A => lbl0_n_19, B => lbl0_n_12, CO => lbl0_n_75, S => lbl0_n_77);
  lbl0_g11070 : INR2XD0BWP7T port map(A1 => lbl0_n_16, B1 => lbl0_n_53, ZN => lbl0_n_71);
  lbl0_g11071 : NR2XD0BWP7T port map(A1 => lbl0_n_53, A2 => lbl0_unsigned_busy_count(0), ZN => lbl0_n_70);
  lbl0_g11072 : INR2D0BWP7T port map(A1 => lbl0_n_57, B1 => memory_ready, ZN => lbl0_n_69);
  lbl0_g11073 : INR2XD0BWP7T port map(A1 => lbl0_n_58, B1 => lbl0_n_53, ZN => lbl0_n_68);
  lbl0_g11074 : INR2D1BWP7T port map(A1 => lbl0_n_50, B1 => lbl0_state(4), ZN => lbl0_n_74);
  lbl0_g11075 : IND2D1BWP7T port map(A1 => lbl0_n_53, B1 => lbl0_counter_busy_counter_state(0), ZN => lbl0_n_72);
  lbl0_g11076 : AOI21D0BWP7T port map(A1 => busy, A2 => lbl0_n_33, B => lbl0_n_32, ZN => lbl0_n_63);
  lbl0_g11077 : OAI211D1BWP7T port map(A1 => lbl0_n_517, A2 => lbl0_n_6, B => lbl0_n_39, C => lbl0_n_56, ZN => FE_PHN78_lbl0_n_62);
  lbl0_g11078 : INR2XD0BWP7T port map(A1 => lbl0_n_38, B1 => lbl0_n_53, ZN => lbl0_n_61);
  lbl0_g11079 : OAI211D1BWP7T port map(A1 => lbl0_n_17, A2 => lbl0_n_5, B => lbl0_n_23, C => lbl0_state(1), ZN => lbl0_n_67);
  lbl0_g11080 : NR4D0BWP7T port map(A1 => lbl0_n_20, A2 => lbl0_mem_com_state(2), A3 => lbl0_mem_com_state(1), A4 => FE_OFN3_rst, ZN => lbl0_n_66);
  lbl0_g11081 : ND2D1BWP7T port map(A1 => lbl0_n_47, A2 => lbl0_state(3), ZN => lbl0_n_65);
  lbl0_g11082 : IND2D1BWP7T port map(A1 => lbl0_n_58, B1 => lbl0_unsigned_busy_count(4), ZN => lbl0_n_64);
  lbl0_g11084 : INVD1BWP7T port map(I => lbl0_n_56, ZN => lbl0_n_57);
  lbl0_g11085 : INR2D1BWP7T port map(A1 => lbl0_n_476, B1 => lbl0_n_30, ZN => lbl0_n_52);
  lbl0_g11086 : OR4D1BWP7T port map(A1 => FE_PHN50_lbl0_unsigned_busy_count_2, A2 => lbl0_unsigned_busy_count(1), A3 => lbl0_n_476, A4 => lbl0_n_477, Z => lbl0_n_51);
  lbl0_g11087 : INR2XD0BWP7T port map(A1 => lbl0_n_40, B1 => lbl0_n_512, ZN => lbl0_n_60);
  lbl0_g11089 : IND2D1BWP7T port map(A1 => lbl0_n_38, B1 => lbl0_unsigned_busy_count(3), ZN => lbl0_n_58);
  lbl0_g11090 : IND3D1BWP7T port map(A1 => lbl0_mem_com_state(1), B1 => FE_PHN82_lbl0_mem_com_state_2, B2 => lbl0_n_18, ZN => lbl0_n_56);
  lbl0_g11091 : IND3D1BWP7T port map(A1 => lbl0_n_14, B1 => lbl0_n_26, B2 => lbl0_n_437, ZN => lbl0_n_55);
  lbl0_g11092 : INR2XD0BWP7T port map(A1 => lbl0_n_33, B1 => lbl0_n_32, ZN => lbl0_n_54);
  lbl0_g11093 : IND2D1BWP7T port map(A1 => lbl0_n_32, B1 => lbl0_counter_busy_counter_state(1), ZN => lbl0_n_53);
  lbl0_g11094 : AOI21D0BWP7T port map(A1 => lbl0_n_28, A2 => lbl0_n_511, B => lbl0_n_509, ZN => lbl0_n_46);
  lbl0_g11095 : AOI22D0BWP7T port map(A1 => lbl0_n_22, A2 => lbl0_state(1), B1 => lbl0_n_5, B2 => lbl0_n_430, ZN => lbl0_n_45);
  lbl0_g11096 : AO21D0BWP7T port map(A1 => lbl0_n_12, A2 => lbl0_n_26, B => lbl0_n_25, Z => lbl0_n_44);
  lbl0_g11097 : MOAI22D0BWP7T port map(A1 => lbl0_n_9, A2 => lbl0_n_10, B1 => lbl0_n_22, B2 => lbl0_n_25, ZN => lbl0_n_43);
  lbl0_g11099 : ND3D0BWP7T port map(A1 => lbl0_n_511, A2 => lbl0_n_27, A3 => start_in, ZN => lbl0_n_41);
  lbl0_g11100 : AN3D0BWP7T port map(A1 => lbl0_n_26, A2 => lbl0_state(1), A3 => lbl0_state(3), Z => lbl0_n_50);
  lbl0_g11101 : ND3D0BWP7T port map(A1 => lbl0_n_427, A2 => lbl0_n_23, A3 => lbl0_state(1), ZN => lbl0_n_49);
  lbl0_g11102 : ND3D0BWP7T port map(A1 => lbl0_n_436, A2 => lbl0_state(1), A3 => lbl0_n_11, ZN => lbl0_n_48);
  lbl0_g11103 : INR3D0BWP7T port map(A1 => lbl0_n_26, B1 => lbl0_state(4), B2 => lbl0_n_8, ZN => lbl0_n_47);
  lbl0_g11104 : AN2D0BWP7T port map(A1 => lbl0_n_15, A2 => lbl0_n_5, Z => lbl0_n_37);
  lbl0_g11105 : IND3D1BWP7T port map(A1 => lbl0_counter_busy_counter_state(1), B1 => lbl0_counter_busy_counter_state(0), B2 => busy, ZN => lbl0_n_36);
  lbl0_g11106 : IND3D0BWP7T port map(A1 => lbl0_state(2), B1 => lbl0_n_13, B2 => lbl0_n_505, ZN => lbl0_n_40);
  lbl0_g11107 : ND2D1BWP7T port map(A1 => lbl0_n_15, A2 => lbl0_mem_com_n_166, ZN => lbl0_n_39);
  lbl0_g11108 : IND2D1BWP7T port map(A1 => lbl0_n_16, B1 => FE_PHN50_lbl0_unsigned_busy_count_2, ZN => lbl0_n_38);
  lbl0_g11109 : OA21D0BWP7T port map(A1 => lbl0_n_504, A2 => lbl0_n_417, B => FE_DBTN4_rst, Z => lbl0_n_31);
  lbl0_g11110 : AOI21D0BWP7T port map(A1 => lbl0_n_477, A2 => lbl0_unsigned_busy_count(0), B => lbl0_unsigned_busy_count(1), ZN => lbl0_n_30);
  lbl0_g11111 : AN3D0BWP7T port map(A1 => lbl0_n_427, A2 => lbl0_n_430, A3 => FE_DBTN4_rst, Z => lbl0_n_35);
  lbl0_g11112 : IND3D1BWP7T port map(A1 => FE_PHN60_lbl0_booster_0, B1 => FE_DBTN4_rst, B2 => lbl0_n_508, ZN => lbl0_n_34);
  lbl0_g11113 : MAOI22D0BWP7T port map(A1 => lbl0_counter_busy_counter_state(1), A2 => lbl0_counter_busy_counter_state(0), B1 => lbl0_counter_busy_counter_state(1), B2 => lbl0_counter_busy_counter_state(0), ZN => lbl0_n_33);
  lbl0_g11114 : OAI21D0BWP7T port map(A1 => lbl0_n_410, A2 => lbl0_n_419, B => FE_DBTN4_rst, ZN => lbl0_n_32);
  lbl0_g11115 : INVD0BWP7T port map(I => lbl0_n_27, ZN => lbl0_n_28);
  lbl0_g11116 : INVD0BWP7T port map(I => lbl0_n_517, ZN => lbl0_n_23);
  lbl0_g11117 : INVD0BWP7T port map(I => lbl0_n_22, ZN => lbl0_n_21);
  lbl0_g11118 : IND2D1BWP7T port map(A1 => lbl0_mem_com_state(0), B1 => lbl0_mem_com_state(3), ZN => lbl0_n_20);
  lbl0_g11119 : NR2XD0BWP7T port map(A1 => lbl0_unsigned_busy_count(5), A2 => lbl0_unsigned_busy_count(6), ZN => lbl0_n_29);
  lbl0_g11120 : NR2D1BWP7T port map(A1 => lbl0_n_428, A2 => lbl0_n_429, ZN => lbl0_n_27);
  lbl0_g11121 : AN2D1BWP7T port map(A1 => player_state_0(0), A2 => player_state_0(1), Z => lbl0_n_19);
  lbl0_g11122 : AN2D1BWP7T port map(A1 => lbl0_state(2), A2 => FE_DBTN4_rst, Z => lbl0_n_26);
  lbl0_g11123 : NR2D1BWP7T port map(A1 => lbl0_n_8, A2 => FE_OFN3_rst, ZN => lbl0_n_25);
  lbl0_g11125 : NR2D1BWP7T port map(A1 => lbl0_n_1952_BAR, A2 => lbl0_state(3), ZN => lbl0_n_22);
  lbl0_g11126 : INVD0BWP7T port map(I => lbl0_n_14, ZN => lbl0_n_13);
  lbl0_g11127 : INVD1BWP7T port map(I => lbl0_n_11, ZN => lbl0_n_10);
  lbl0_g11128 : NR2XD0BWP7T port map(A1 => lbl0_n_511, A2 => lbl0_n_426, ZN => lbl0_n_9);
  lbl0_g11129 : NR2XD0BWP7T port map(A1 => lbl0_mem_com_state(3), A2 => FE_OFN3_rst, ZN => lbl0_n_18);
  lbl0_g11130 : INR2D1BWP7T port map(A1 => lbl0_booster_1, B1 => lbl0_state(0), ZN => lbl0_n_17);
  lbl0_g11131 : ND2D1BWP7T port map(A1 => lbl0_unsigned_busy_count(1), A2 => lbl0_unsigned_busy_count(0), ZN => lbl0_n_16);
  lbl0_g11132 : AN2D1BWP7T port map(A1 => lbl0_n_513, A2 => FE_DBTN4_rst, Z => lbl0_n_15);
  lbl0_g11133 : ND2D1BWP7T port map(A1 => lbl0_n_8, A2 => lbl0_n_4, ZN => lbl0_n_14);
  lbl0_g11134 : AN2D1BWP7T port map(A1 => player_state_1(0), A2 => player_state_1(1), Z => lbl0_n_12);
  lbl0_g11135 : NR2D0BWP7T port map(A1 => FE_OFN3_rst, A2 => start_in, ZN => lbl0_n_11);
  lbl0_g11139 : INVD0BWP7T port map(I => lbl0_mem_com_n_166, ZN => lbl0_n_6);
  lbl0_g11140 : INVD1BWP7T port map(I => lbl0_n_427, ZN => lbl0_n_5);
  lbl0_g14949 : IND3D1BWP7T port map(A1 => lbl0_n_103, B1 => lbl0_n_510, B2 => FE_DBTN4_rst, ZN => lbl0_n_1);
  lbl0_g11145 : IND3D1BWP7T port map(A1 => lbl0_n_60, B1 => FE_DBTN4_rst, B2 => start_in, ZN => lbl0_n_0);
  lbl0_g14950 : OR2D1BWP7T port map(A1 => lbl0_n_11, A2 => lbl0_n_25, Z => lbl0_n_515);
  lbl0_mem_com_state_reg_0 : DFD1BWP7T port map(CP => CTS_12, D => lbl0_n_122, Q => lbl0_mem_com_state(0), QN => lbl0_n_160);
  lbl0_mem_com_state_reg_1 : DFD1BWP7T port map(CP => CTS_12, D => lbl0_n_110, Q => lbl0_mem_com_state(1), QN => lbl0_n_157);
  lbl0_state_reg_4 : DFD1BWP7T port map(CP => CTS_11, D => lbl0_n_133, Q => lbl0_state(4), QN => lbl0_n_156);
  lbl0_mem_com_state_reg_2 : DFD1BWP7T port map(CP => CTS_12, D => lbl0_n_62, Q => lbl0_mem_com_state(2), QN => lbl0_n_152);
  lbl0_state_reg_3 : DFD1BWP7T port map(CP => CTS_11, D => lbl0_n_129, Q => lbl0_state(3), QN => lbl0_n_147);
  lbl0_state_reg_0 : DFD1BWP7T port map(CP => CTS_12, D => lbl0_n_131, Q => lbl0_state(0), QN => lbl0_n_8);
  lbl0_counter_unsigned_busy_count_reg_0 : DFD1BWP7T port map(CP => CTS_11, D => lbl0_n_94, Q => FE_PHN47_lbl0_unsigned_busy_count_0, QN => lbl0_n_7);
  lbl0_state_reg_1 : DFD1BWP7T port map(CP => CTS_11, D => lbl0_n_132, Q => lbl0_state(1), QN => lbl0_n_4);
  lbl0_g14967 : INR4D0BWP7T port map(A1 => lbl0_n_15, B1 => lbl0_n_194, B2 => lbl0_mem_com_state(2), B3 => lbl0_mem_com_state(1), ZN => lbl0_n_516);
  lbl0_g14968 : IND3D1BWP7T port map(A1 => lbl0_state(2), B1 => lbl0_n_437, B2 => FE_DBTN4_rst, ZN => lbl0_n_517);
  lbl0_reg_pos0_q_reg_2 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_0(2), E => lbl0_e_position_0, Q => position_0(2));
  lbl0_reg_pos0_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_0(1), E => lbl0_e_position_0, Q => position_0(1));
  lbl0_reg_pos0_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_n_411, E => lbl0_e_position_0, Q => position_0(0));
  lbl0_reg_pos0_q_reg_7 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_0(7), E => lbl0_e_position_0, Q => position_0(7));
  lbl0_reg_pos0_q_reg_8 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_0(8), E => lbl0_e_position_0, Q => position_0(8));
  lbl0_reg_pos0_q_reg_4 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_n_412, E => lbl0_e_position_0, Q => position_0(4));
  lbl0_reg_pos0_q_reg_3 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_0(3), E => lbl0_e_position_0, Q => position_0(3));
  lbl0_reg_pos0_q_reg_9 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_n_414, E => lbl0_e_position_0, Q => position_0(9));
  lbl0_reg_pos0_q_reg_5 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_n_413, E => lbl0_e_position_0, Q => position_0(5));
  lbl0_reg_pos0_q_reg_6 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_0(6), E => lbl0_e_position_0, Q => position_0(6));
  lbl0_reg_n_layer_1_q_reg : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_n_473, E => lbl0_n_506, Q => lbl0_next_layer_1);
  lbl0_reg_booster_sync_q_reg : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_booster_sync, E => lbl0_n_432, Q => lbl0_booster_sync);
  lbl0_reg_pos1_q_reg_2 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_1(2), E => lbl0_e_position_1, Q => position_1(2));
  lbl0_reg_pos1_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_1(1), E => lbl0_e_position_1, Q => position_1(1));
  lbl0_reg_pos1_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_1(0), E => lbl0_e_position_1, Q => position_1(0));
  lbl0_reg_pos1_q_reg_7 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_1(7), E => lbl0_e_position_1, Q => position_1(7));
  lbl0_reg_pos1_q_reg_8 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_1(8), E => lbl0_e_position_1, Q => position_1(8));
  lbl0_reg_pos1_q_reg_4 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_1(4), E => lbl0_e_position_1, Q => position_1(4));
  lbl0_reg_pos1_q_reg_3 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_1(3), E => lbl0_e_position_1, Q => position_1(3));
  lbl0_reg_pos1_q_reg_9 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_1(9), E => lbl0_e_position_1, Q => position_1(9));
  lbl0_reg_pos1_q_reg_5 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_1(5), E => lbl0_e_position_1, Q => position_1(5));
  lbl0_reg_pos1_q_reg_6 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_position_1(6), E => lbl0_e_position_1, Q => position_1(6));
  lbl0_reg_booster_0_q_reg : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_booster_0, E => lbl0_n_432, Q => lbl0_booster_0);
  lbl0_reg_border_0_q_reg : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_n_472, E => lbl0_n_507, Q => lbl0_border_0);
  lbl0_reg_booster_1_q_reg : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_booster_1, E => lbl0_n_432, Q => lbl0_booster_1);
  lbl0_reg_border_1_q_reg : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_n_471, E => lbl0_n_506, Q => lbl0_border_1);
  lbl0_reg_dir_0_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_direction_0(0), E => lbl0_n_433, Q => direction_0(0));
  lbl0_reg_dir_0_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_direction_0(1), E => lbl0_n_433, Q => direction_0(1));
  lbl0_reg_p_state_0_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_n_421, E => lbl0_n_416, Q => player_state_0(0));
  lbl0_reg_p_state_0_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_n_422, E => lbl0_n_416, Q => player_state_0(1));
  lbl0_reg_dir_1_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_direction_1(0), E => lbl0_n_433, Q => direction_1(0));
  lbl0_reg_dir_1_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_direction_1(1), E => lbl0_n_433, Q => direction_1(1));
  lbl0_reg_speed_select_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_speed_select(0), E => lbl0_n_512, Q => lbl0_n_477);
  lbl0_reg_speed_select_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_speed_select(1), E => lbl0_n_512, Q => lbl0_n_476);
  lbl0_reg_p_state_1_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_n_420, E => lbl0_n_415, Q => player_state_1(0));
  lbl0_reg_p_state_1_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_n_422, E => lbl0_n_415, Q => player_state_1(1));
  lbl0_reg_n_dir_0_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_next_direction_0(0), E => lbl0_n_425, Q => lbl0_next_direction_0(0));
  lbl0_reg_n_dir_0_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_next_direction_0(1), E => lbl0_n_425, Q => lbl0_next_direction_0(1));
  lbl0_reg_layer_0_q_reg : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_layer_0, E => lbl0_e_position_0, Q => position_0(10));
  lbl0_reg_n_dir_1_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_next_direction_1(0), E => lbl0_n_424, Q => lbl0_next_direction_1(0));
  lbl0_reg_n_dir_1_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_next_direction_1(1), E => lbl0_n_424, Q => lbl0_next_direction_1(1));
  lbl0_reg_layer_1_q_reg : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_11, D => lbl0_d_layer_1, E => lbl0_e_position_1, Q => position_1(10));
  lbl0_reg_map_select_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_map_select(0), E => lbl0_n_512, Q => map_selected(0));
  lbl0_reg_map_select_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_map_select(1), E => lbl0_n_512, Q => map_selected(1));
  lbl0_reg_r_mem_0_q_reg_3 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_read_data_reg(3), E => lbl0_n_430, Q => lbl0_read_data_reg(3));
  lbl0_reg_r_mem_0_q_reg_2 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_read_data_reg(2), E => lbl0_n_430, Q => lbl0_read_data_reg(2));
  lbl0_reg_r_mem_0_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_read_data_reg(0), E => lbl0_n_430, Q => lbl0_read_data_reg(0));
  lbl0_reg_r_mem_0_q_reg_4 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_read_data_reg(4), E => lbl0_n_430, Q => lbl0_read_data_reg(4));
  lbl0_reg_r_mem_0_q_reg_6 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_read_data_reg(6), E => lbl0_n_430, Q => lbl0_read_data_reg(6));
  lbl0_reg_r_mem_0_q_reg_5 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_read_data_reg(5), E => lbl0_n_430, Q => lbl0_read_data_reg(5));
  lbl0_reg_r_mem_0_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_read_data_reg(1), E => lbl0_n_430, Q => lbl0_read_data_reg(1));
  lbl0_reg_r_mem_0_q_reg_7 : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_d_read_data_reg(7), E => lbl0_n_430, Q => lbl0_read_data_reg(7));
  lbl1_g14 : INVD1BWP7T port map(I => memory_ready, ZN => lbl1_n_1);
  lbl1_g19 : CKAN2D1BWP7T port map(A1 => lbl1_ready_rw, A2 => lbl1_ready_clr, Z => memory_ready);
  lbl1_g22 : OR3D4BWP7T port map(A1 => lbl1_x_incr3, A2 => lbl1_x_incr2, A3 => lbl1_x_incr1, Z => x_increment_out);
  lbl1_g23 : OR3D4BWP7T port map(A1 => lbl1_y_incr3, A2 => lbl1_y_incr2, A3 => lbl1_y_incr1, Z => y_increment_out);
  lbl1_g24 : CKAN2D8BWP7T port map(A1 => lbl1_we_clr, A2 => lbl1_we_rw, Z => write_enable_out);
  lbl1_g13 : OR2D1BWP7T port map(A1 => lbl1_me_rw, A2 => lbl1_me_clr, Z => FE_OFN5_memory_enable_out);
  lbl1_g27 : OR4D4BWP7T port map(A1 => FE_OFN3_rst, A2 => lbl1_clr_rst, A3 => lbl1_rw_rst, A4 => reset_vga_mem, Z => memory_reset_out);
  lbl1_cy_count_reg_4 : DFCNQD1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => y_increment_out, D => lbl1_cy_n_8, Q => y_address(4));
  lbl1_cy_g82 : MOAI22D0BWP7T port map(A1 => lbl1_cy_n_6, A2 => y_address(4), B1 => lbl1_cy_n_6, B2 => y_address(4), ZN => lbl1_cy_n_8);
  lbl1_cy_count_reg_3 : DFCNQD1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => y_increment_out, D => lbl1_cy_n_7, Q => y_address(3));
  lbl1_cy_g84 : MOAI22D0BWP7T port map(A1 => lbl1_cy_n_4, A2 => y_address(3), B1 => lbl1_cy_n_4, B2 => y_address(3), ZN => lbl1_cy_n_7);
  lbl1_cy_count_reg_2 : DFCNQD1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => y_increment_out, D => lbl1_cy_n_5, Q => y_address(2));
  lbl1_cy_g86 : IND2D0BWP7T port map(A1 => lbl1_cy_n_4, B1 => y_address(3), ZN => lbl1_cy_n_6);
  lbl1_cy_g87 : MOAI22D0BWP7T port map(A1 => lbl1_cy_n_3, A2 => y_address(2), B1 => lbl1_cy_n_3, B2 => y_address(2), ZN => lbl1_cy_n_5);
  lbl1_cy_g89 : IND2D0BWP7T port map(A1 => lbl1_cy_n_3, B1 => y_address(2), ZN => lbl1_cy_n_4);
  lbl1_cy_g91 : ND2D0BWP7T port map(A1 => y_address(0), A2 => y_address(1), ZN => lbl1_cy_n_3);
  lbl1_cy_count_reg_1 : EDFCND1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => y_increment_out, D => lbl1_cy_n_2, E => y_address(0), Q => y_address(1), QN => lbl1_cy_n_2);
  lbl1_cy_count_reg_0 : DFCND1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => y_increment_out, D => lbl1_cy_n_0, Q => y_address(0), QN => lbl1_cy_n_0);
  lbl1_cm_g544 : AO221D0BWP7T port map(A1 => lbl1_cm_n_37, A2 => lbl1_cm_n_28, B1 => lbl1_cm_n_29, B2 => lbl1_cm_state(3), C => lbl1_x_incr3, Z => lbl1_we_clr);
  lbl1_cm_g545 : AO31D1BWP7T port map(A1 => lbl1_cm_n_28, A2 => lbl1_cm_n_27, A3 => lbl1_cm_state(0), B => lbl1_cm_state(4), Z => lbl1_clr_rst);
  lbl1_cm_g546 : INR4D0BWP7T port map(A1 => lbl1_cm_n_28, B1 => lbl1_cm_state(1), B2 => lbl1_cm_state(0), B3 => lbl1_cm_state(4), ZN => lbl1_ready_clr);
  lbl1_cm_g547 : AN2D0BWP7T port map(A1 => lbl1_x_incr3, A2 => lbl1_cm_state(1), Z => lbl1_y_incr3);
  lbl1_cm_g548 : CKND1BWP7T port map(I => lbl1_cm_n_37, ZN => lbl1_cm_n_29);
  lbl1_cm_g549 : NR2XD0BWP7T port map(A1 => lbl1_cm_n_27, A2 => lbl1_cm_state(2), ZN => lbl1_me_clr);
  lbl1_cm_g550 : ND2D1BWP7T port map(A1 => lbl1_cm_state(0), A2 => lbl1_cm_state(1), ZN => lbl1_cm_n_37);
  lbl1_cm_g551 : IND2D1BWP7T port map(A1 => lbl1_cm_state(3), B1 => lbl1_cm_state(0), ZN => lbl1_cm_n_32);
  lbl1_cm_g552 : CKAN2D1BWP7T port map(A1 => lbl1_cm_state(2), A2 => lbl1_cm_state(3), Z => lbl1_x_incr3);
  lbl1_cm_g553 : NR2XD0BWP7T port map(A1 => lbl1_cm_state(2), A2 => lbl1_cm_state(3), ZN => lbl1_cm_n_28);
  lbl1_cm_state_reg_2 : DFQD1BWP7T port map(CP => CTS_12, D => FE_PHN43_lbl1_cm_n_25, Q => lbl1_cm_state(2));
  lbl1_cm_state_reg_0 : DFQD1BWP7T port map(CP => CTS_12, D => FE_PHN72_lbl1_cm_n_24, Q => lbl1_cm_state(0));
  lbl1_cm_g809 : OAI211D1BWP7T port map(A1 => lbl1_cm_n_10, A2 => lbl1_cm_n_13, B => lbl1_cm_n_15, C => lbl1_cm_n_22, ZN => lbl1_cm_n_26);
  lbl1_cm_state_reg_4 : DFKCNQD1BWP7T port map(CN => lbl1_cm_n_20, CP => CTS_12, D => lbl1_cm_n_17, Q => lbl1_cm_state(4));
  lbl1_cm_g811 : OAI211D1BWP7T port map(A1 => lbl1_cm_n_9, A2 => lbl1_cm_n_13, B => lbl1_cm_n_14, C => lbl1_cm_n_22, ZN => lbl1_cm_n_25);
  lbl1_cm_g812 : MOAI22D0BWP7T port map(A1 => lbl1_cm_n_11, A2 => FE_OFN3_rst, B1 => lbl1_cm_n_5, B2 => lbl1_cm_n_52, ZN => lbl1_cm_n_24);
  lbl1_cm_g813 : OAI32D1BWP7T port map(A1 => lbl1_cm_n_8, A2 => lbl1_cm_n_12, A3 => lbl1_cm_n_4, B1 => lbl1_cm_n_18, B2 => lbl1_cm_n_21, ZN => FE_PHN48_lbl1_cm_n_23);
  lbl1_cm_g814 : IND2D1BWP7T port map(A1 => lbl1_cm_n_20, B1 => lbl1_cm_n_17, ZN => lbl1_cm_n_22);
  lbl1_cm_g815 : ND2D1BWP7T port map(A1 => lbl1_cm_n_17, A2 => lbl1_cm_n_16, ZN => lbl1_cm_n_21);
  lbl1_cm_g817 : NR2D0BWP7T port map(A1 => lbl1_cm_n_18, A2 => lbl1_cm_n_16, ZN => lbl1_cm_n_20);
  lbl1_cm_g818 : IND4D0BWP7T port map(A1 => lbl1_cm_n_6, B1 => x_address(3), B2 => x_address(0), B3 => x_address(1), ZN => lbl1_cm_n_18);
  lbl1_cm_g819 : INR2XD0BWP7T port map(A1 => lbl1_cm_n_12, B1 => FE_OFN3_rst, ZN => lbl1_cm_n_17);
  lbl1_cm_g820 : IND4D0BWP7T port map(A1 => lbl1_cm_state(2), B1 => lbl1_cm_state(3), B2 => lbl1_cm_n_37, B3 => lbl1_cm_n_5, ZN => lbl1_cm_n_15);
  lbl1_cm_g821 : IND3D1BWP7T port map(A1 => lbl1_cm_state(2), B1 => lbl1_cm_n_7, B2 => lbl1_cm_n_5, ZN => lbl1_cm_n_14);
  lbl1_cm_g822 : IND4D0BWP7T port map(A1 => lbl1_cm_n_3, B1 => y_address(2), B2 => y_address(1), B3 => y_address(4), ZN => lbl1_cm_n_16);
  lbl1_cm_g823 : IND3D1BWP7T port map(A1 => lbl1_n_1, B1 => clear_memory, B2 => lbl1_ready_clr, ZN => lbl1_cm_n_11);
  lbl1_cm_g824 : ND2D1BWP7T port map(A1 => lbl1_cm_n_5, A2 => lbl1_cm_state(2), ZN => lbl1_cm_n_13);
  lbl1_cm_g825 : NR3D0BWP7T port map(A1 => lbl1_cm_n_37, A2 => lbl1_cm_n_2, A3 => lbl1_cm_state(2), ZN => lbl1_cm_n_12);
  lbl1_cm_g826 : IAO21D0BWP7T port map(A1 => lbl1_cm_n_2, A2 => lbl1_cm_state(0), B => lbl1_cm_n_7, ZN => lbl1_cm_n_10);
  lbl1_cm_g827 : OA21D0BWP7T port map(A1 => lbl1_cm_state(1), A2 => lbl1_cm_state(3), B => lbl1_cm_state(0), Z => lbl1_cm_n_9);
  lbl1_cm_g828 : MUX2ND0BWP7T port map(I0 => lbl1_cm_state(0), I1 => lbl1_cm_n_32, S => lbl1_cm_state(1), ZN => lbl1_cm_n_8);
  lbl1_cm_g829 : ND2D0BWP7T port map(A1 => x_address(2), A2 => x_address(4), ZN => lbl1_cm_n_6);
  lbl1_cm_g830 : NR2D1BWP7T port map(A1 => lbl1_cm_n_37, A2 => lbl1_cm_state(3), ZN => lbl1_cm_n_7);
  lbl1_cm_g831 : INVD0BWP7T port map(I => lbl1_cm_n_5, ZN => lbl1_cm_n_4);
  lbl1_cm_g832 : ND2D0BWP7T port map(A1 => y_address(0), A2 => y_address(3), ZN => lbl1_cm_n_3);
  lbl1_cm_g833 : NR2XD0BWP7T port map(A1 => lbl1_ready_clr, A2 => FE_OFN3_rst, ZN => lbl1_cm_n_5);
  lbl1_cm_g2 : NR2D1BWP7T port map(A1 => lbl1_cm_state(0), A2 => lbl1_cm_state(4), ZN => lbl1_cm_n_52);
  lbl1_cm_state_reg_1 : DFD1BWP7T port map(CP => CTS_12, D => lbl1_cm_n_23, Q => lbl1_cm_state(1), QN => lbl1_cm_n_27);
  lbl1_cm_state_reg_3 : DFD1BWP7T port map(CP => CTS_12, D => FE_PHN40_lbl1_cm_n_26, Q => lbl1_cm_state(3), QN => lbl1_cm_n_2);
  lbl1_cex_g177 : OR2D1BWP7T port map(A1 => lbl1_cex_n_9, A2 => lbl1_cex_n_8, Z => lbl1_x_incr2);
  lbl1_cex_g178 : INR2D1BWP7T port map(A1 => lbl1_cex_state(1), B1 => lbl1_cex_state(0), ZN => lbl1_cex_n_8);
  lbl1_cex_g179 : INR2D1BWP7T port map(A1 => lbl1_cex_state(0), B1 => lbl1_cex_state(1), ZN => lbl1_cex_n_9);
  lbl1_cex_state_reg_0 : DFQD1BWP7T port map(CP => CTS_11, D => lbl1_cex_n_7, Q => lbl1_cex_state(0));
  lbl1_cex_g169 : NR2XD0BWP7T port map(A1 => FE_PHN74_lbl1_cex_n_6, A2 => FE_OFN3_rst, ZN => lbl1_cex_n_7);
  lbl1_cex_g171 : AOI21D0BWP7T port map(A1 => x_increment, A2 => lbl1_cex_n_4, B => FE_PHN37_lbl1_cex_n_8, ZN => lbl1_cex_n_6);
  lbl1_cex_g172 : NR2XD0BWP7T port map(A1 => FE_PHN68_lbl1_cex_n_3, A2 => FE_OFN3_rst, ZN => lbl1_cex_n_5);
  lbl1_cex_g173 : AOI21D0BWP7T port map(A1 => lbl1_n_1, A2 => lbl1_cex_n_2, B => lbl1_cex_n_9, ZN => lbl1_cex_n_4);
  lbl1_cex_g174 : AOI21D0BWP7T port map(A1 => x_increment, A2 => lbl1_cex_state(0), B => lbl1_x_incr2, ZN => lbl1_cex_n_3);
  lbl1_cex_state_reg_1 : DFD1BWP7T port map(CP => CTS_11, D => lbl1_cex_n_5, Q => lbl1_cex_state(1), QN => lbl1_cex_n_2);
  lbl1_rw_g1135 : OAI21D0BWP7T port map(A1 => lbl1_rw_n_81, A2 => lbl1_rw_n_100, B => lbl1_rw_n_87, ZN => lbl1_me_rw);
  lbl1_rw_g1136 : NR3D0BWP7T port map(A1 => lbl1_rw_n_82, A2 => lbl1_rw_n_90, A3 => lbl1_rw_state(4), ZN => lbl1_rw_rst);
  lbl1_rw_g1137 : NR3D0BWP7T port map(A1 => lbl1_rw_n_82, A2 => lbl1_rw_state(4), A3 => lbl1_rw_state(0), ZN => lbl1_ready_rw);
  lbl1_rw_g1138 : OAI221D0BWP7T port map(A1 => lbl1_rw_n_77, A2 => lbl1_rw_n_83, B1 => lbl1_rw_n_88, B2 => lbl1_rw_n_84, C => lbl1_rw_n_80, ZN => lbl1_y_incr1);
  lbl1_rw_g1139 : OAI221D0BWP7T port map(A1 => lbl1_rw_n_99, A2 => lbl1_rw_state(4), B1 => lbl1_rw_state(1), B2 => lbl1_rw_n_83, C => lbl1_rw_n_80, ZN => lbl1_x_incr1);
  lbl1_rw_g1140 : MOAI22D0BWP7T port map(A1 => lbl1_rw_n_79, A2 => lbl1_rw_n_90, B1 => lbl1_rw_n_100, B2 => lbl1_rw_n_87, ZN => lbl1_we_rw);
  lbl1_rw_g1141 : IND3D1BWP7T port map(A1 => lbl1_rw_n_77, B1 => lbl1_rw_n_89, B2 => lbl1_rw_n_87, ZN => lbl1_rw_n_82);
  lbl1_rw_g1142 : OAI21D2BWP7T port map(A1 => lbl1_rw_n_83, A2 => lbl1_rw_n_78, B => lbl1_rw_n_80, ZN => w_increment_out);
  lbl1_rw_g1143 : IAO21D0BWP7T port map(A1 => lbl1_rw_n_99, A2 => lbl1_rw_n_90, B => lbl1_rw_n_97, ZN => lbl1_rw_n_81);
  lbl1_rw_g1144 : NR2XD0BWP7T port map(A1 => lbl1_rw_n_86, A2 => lbl1_rw_n_88, ZN => lbl1_rw_n_97);
  lbl1_rw_g1145 : AN2D0BWP7T port map(A1 => lbl1_rw_n_99, A2 => lbl1_rw_n_87, Z => lbl1_rw_n_79);
  lbl1_rw_g1146 : IND2D1BWP7T port map(A1 => lbl1_rw_n_85, B1 => lbl1_rw_n_78, ZN => lbl1_rw_n_80);
  lbl1_rw_g1147 : CKND2D1BWP7T port map(A1 => lbl1_rw_n_89, A2 => lbl1_rw_state(4), ZN => lbl1_rw_n_85);
  lbl1_rw_g1148 : IND2D1BWP7T port map(A1 => lbl1_rw_state(4), B1 => lbl1_rw_state(3), ZN => lbl1_rw_n_83);
  lbl1_rw_g1149 : ND2D1BWP7T port map(A1 => lbl1_rw_n_88, A2 => lbl1_rw_state(2), ZN => lbl1_rw_n_99);
  lbl1_rw_g1150 : INVD0BWP7T port map(I => lbl1_rw_n_78, ZN => lbl1_rw_n_77);
  lbl1_rw_g1151 : ND2D1BWP7T port map(A1 => lbl1_rw_n_90, A2 => lbl1_rw_state(2), ZN => lbl1_rw_n_86);
  lbl1_rw_g1152 : IND2D1BWP7T port map(A1 => lbl1_rw_state(4), B1 => lbl1_rw_state(2), ZN => lbl1_rw_n_84);
  lbl1_rw_g1153 : CKND2D1BWP7T port map(A1 => lbl1_rw_state(4), A2 => lbl1_rw_state(3), ZN => lbl1_rw_n_100);
  lbl1_rw_g1154 : NR2XD0BWP7T port map(A1 => lbl1_rw_state(2), A2 => lbl1_rw_state(1), ZN => lbl1_rw_n_78);
  lbl1_rw_state_reg_2 : DFQD1BWP7T port map(CP => CTS_12, D => lbl1_rw_n_75, Q => lbl1_rw_state(2));
  lbl1_rw_state_reg_4 : DFQD1BWP7T port map(CP => CTS_12, D => lbl1_rw_n_73, Q => lbl1_rw_state(4));
  lbl1_rw_g2250 : ND2D1BWP7T port map(A1 => lbl1_rw_n_72, A2 => lbl1_rw_n_58, ZN => lbl1_rw_n_76);
  lbl1_rw_g2251 : OR4D1BWP7T port map(A1 => lbl1_rw_n_64, A2 => lbl1_rw_n_63, A3 => lbl1_rw_n_68, A4 => lbl1_rw_n_62, Z => lbl1_rw_n_75);
  lbl1_rw_g2252 : ND3D0BWP7T port map(A1 => lbl1_rw_n_66, A2 => lbl1_rw_n_59, A3 => lbl1_rw_n_52, ZN => lbl1_rw_n_74);
  lbl1_rw_g2254 : OR3D1BWP7T port map(A1 => lbl1_rw_n_67, A2 => lbl1_rw_n_69, A3 => FE_PHN79_lbl1_rw_n_0, Z => lbl1_rw_n_73);
  lbl1_rw_g2255 : AOI211XD0BWP7T port map(A1 => lbl1_rw_n_64, A2 => lbl1_rw_n_41, B => lbl1_rw_n_65, C => lbl1_rw_n_61, ZN => lbl1_rw_n_72);
  lbl1_rw_g2256 : OAI211D1BWP7T port map(A1 => FE_OFN3_rst, A2 => lbl1_rw_n_28, B => lbl1_rw_n_56, C => lbl1_rw_n_70, ZN => lbl1_rw_n_71);
  lbl1_rw_g2257 : INVD0BWP7T port map(I => lbl1_rw_n_69, ZN => lbl1_rw_n_70);
  lbl1_rw_g2258 : OAI221D0BWP7T port map(A1 => lbl1_rw_n_52, A2 => lbl1_rw_n_39, B1 => lbl1_rw_n_38, B2 => lbl1_rw_n_49, C => lbl1_rw_n_45, ZN => lbl1_rw_n_68);
  lbl1_rw_g2259 : OAI22D0BWP7T port map(A1 => lbl1_rw_n_58, A2 => lbl1_rw_n_41, B1 => lbl1_rw_n_52, B2 => lbl1_rw_n_38, ZN => lbl1_rw_n_69);
  lbl1_rw_g2261 : OAI211D1BWP7T port map(A1 => lbl1_rw_n_40, A2 => lbl1_rw_n_57, B => lbl1_rw_n_55, C => lbl1_rw_n_46, ZN => lbl1_rw_n_67);
  lbl1_rw_g2262 : MAOI22D0BWP7T port map(A1 => lbl1_rw_n_43, A2 => FE_PHN55_lbl1_rw_n_29, B1 => lbl1_rw_n_58, B2 => lbl1_rw_n_40, ZN => lbl1_rw_n_66);
  lbl1_rw_g2263 : OAI22D0BWP7T port map(A1 => lbl1_rw_n_57, A2 => lbl1_rw_n_41, B1 => lbl1_rw_n_47, B2 => lbl1_rw_n_4, ZN => lbl1_rw_n_65);
  lbl1_rw_g2264 : NR2D0BWP7T port map(A1 => lbl1_rw_n_58, A2 => lbl1_rw_n_41, ZN => lbl1_rw_n_63);
  lbl1_rw_g2265 : IOA21D1BWP7T port map(A1 => lbl1_rw_n_53, A2 => lbl1_rw_n_39, B => lbl1_rw_n_59, ZN => lbl1_rw_n_64);
  lbl1_rw_g2266 : OAI22D0BWP7T port map(A1 => lbl1_rw_n_48, A2 => lbl1_rw_n_88, B1 => lbl1_rw_n_51, B2 => lbl1_rw_n_84, ZN => lbl1_rw_n_62);
  lbl1_rw_g2267 : OAI22D0BWP7T port map(A1 => lbl1_rw_n_49, A2 => lbl1_rw_n_39, B1 => lbl1_rw_n_51, B2 => lbl1_rw_n_83, ZN => lbl1_rw_n_61);
  lbl1_rw_g2268 : OAI22D0BWP7T port map(A1 => lbl1_rw_n_47, A2 => lbl1_rw_n_5, B1 => lbl1_rw_n_51, B2 => lbl1_rw_n_87, ZN => lbl1_rw_n_60);
  lbl1_rw_g2269 : CKND2D1BWP7T port map(A1 => lbl1_rw_n_54, A2 => lbl1_rw_n_38, ZN => lbl1_rw_n_59);
  lbl1_rw_g2270 : ND2D1BWP7T port map(A1 => lbl1_rw_n_54, A2 => lbl1_rw_n_39, ZN => lbl1_rw_n_58);
  lbl1_rw_g2271 : OAI21D0BWP7T port map(A1 => lbl1_rw_n_99, A2 => lbl1_rw_n_100, B => lbl1_rw_n_50, ZN => lbl1_rw_n_56);
  lbl1_rw_g2272 : AO21D0BWP7T port map(A1 => lbl1_rw_n_88, A2 => lbl1_rw_state(2), B => lbl1_rw_n_47, Z => lbl1_rw_n_55);
  lbl1_rw_g2273 : CKND2D1BWP7T port map(A1 => lbl1_rw_n_53, A2 => lbl1_rw_n_38, ZN => lbl1_rw_n_57);
  lbl1_rw_g2274 : INVD0BWP7T port map(I => lbl1_rw_n_51, ZN => lbl1_rw_n_50);
  lbl1_rw_g2275 : NR2XD0BWP7T port map(A1 => lbl1_rw_n_44, A2 => lbl1_rw_n_37, ZN => lbl1_rw_n_54);
  lbl1_rw_g2276 : NR2D1BWP7T port map(A1 => lbl1_rw_n_44, A2 => lbl1_rw_n_36, ZN => lbl1_rw_n_53);
  lbl1_rw_g2277 : ND2D1BWP7T port map(A1 => lbl1_rw_n_42, A2 => lbl1_rw_n_36, ZN => lbl1_rw_n_52);
  lbl1_rw_g2278 : IND2D1BWP7T port map(A1 => lbl1_rw_state(0), B1 => lbl1_rw_n_43, ZN => lbl1_rw_n_51);
  lbl1_rw_g2279 : INVD0BWP7T port map(I => lbl1_rw_n_0, ZN => lbl1_rw_n_48);
  lbl1_rw_g2280 : OAI21D0BWP7T port map(A1 => lbl1_rw_n_26, A2 => lbl1_rw_n_27, B => lbl1_rw_n_43, ZN => lbl1_rw_n_46);
  lbl1_rw_g2281 : OAI21D0BWP7T port map(A1 => lbl1_rw_n_30, A2 => lbl1_rw_n_97, B => lbl1_rw_n_43, ZN => lbl1_rw_n_45);
  lbl1_rw_g2282 : CKND2D1BWP7T port map(A1 => lbl1_rw_n_42, A2 => lbl1_rw_n_37, ZN => lbl1_rw_n_49);
  lbl1_rw_g2284 : IND2D1BWP7T port map(A1 => lbl1_rw_n_100, B1 => lbl1_rw_n_43, ZN => lbl1_rw_n_47);
  lbl1_rw_g2286 : IND3D1BWP7T port map(A1 => FE_OFN3_rst, B1 => write_enable, B2 => lbl1_rw_n_35, ZN => lbl1_rw_n_44);
  lbl1_rw_g2287 : NR3D0BWP7T port map(A1 => lbl1_ready_rw, A2 => lbl1_rw_n_35, A3 => FE_OFN3_rst, ZN => lbl1_rw_n_43);
  lbl1_rw_g2288 : INVD0BWP7T port map(I => lbl1_rw_n_41, ZN => lbl1_rw_n_40);
  lbl1_rw_g2289 : INR3D0BWP7T port map(A1 => lbl1_rw_n_35, B1 => FE_OFN3_rst, B2 => write_enable, ZN => lbl1_rw_n_42);
  lbl1_rw_g2290 : ND4D0BWP7T port map(A1 => lbl1_rw_n_34, A2 => lbl1_rw_n_31, A3 => lbl1_rw_n_9, A4 => lbl1_rw_n_8, ZN => lbl1_rw_n_41);
  lbl1_rw_g2291 : INVD1BWP7T port map(I => lbl1_rw_n_39, ZN => lbl1_rw_n_38);
  lbl1_rw_g2292 : NR4D0BWP7T port map(A1 => lbl1_rw_n_33, A2 => lbl1_rw_n_17, A3 => lbl1_rw_n_13, A4 => lbl1_rw_n_19, ZN => lbl1_rw_n_39);
  lbl1_rw_g2293 : INVD1BWP7T port map(I => lbl1_rw_n_37, ZN => lbl1_rw_n_36);
  lbl1_rw_g2294 : ND4D0BWP7T port map(A1 => lbl1_rw_n_32, A2 => lbl1_rw_n_10, A3 => lbl1_rw_n_12, A4 => lbl1_rw_n_11, ZN => lbl1_rw_n_37);
  lbl1_rw_g2295 : NR4D0BWP7T port map(A1 => lbl1_rw_n_3, A2 => lbl1_rw_n_88, A3 => lbl1_rw_n_90, A4 => lbl1_rw_state(2), ZN => lbl1_rw_n_35);
  lbl1_rw_g2296 : NR4D0BWP7T port map(A1 => lbl1_rw_n_20, A2 => lbl1_rw_n_21, A3 => lbl1_rw_n_22, A4 => lbl1_rw_n_23, ZN => lbl1_rw_n_34);
  lbl1_rw_g2297 : ND2D1BWP7T port map(A1 => lbl1_rw_n_15, A2 => lbl1_rw_n_16, ZN => lbl1_rw_n_33);
  lbl1_rw_g2298 : NR2XD0BWP7T port map(A1 => lbl1_rw_n_18, A2 => lbl1_rw_n_14, ZN => lbl1_rw_n_32);
  lbl1_rw_g2299 : NR2XD0BWP7T port map(A1 => lbl1_rw_n_25, A2 => lbl1_rw_n_24, ZN => lbl1_rw_n_31);
  lbl1_rw_g2300 : AOI21D0BWP7T port map(A1 => lbl1_rw_n_85, A2 => lbl1_rw_n_7, B => lbl1_rw_n_99, ZN => lbl1_rw_n_30);
  lbl1_rw_g2301 : OAI32D1BWP7T port map(A1 => lbl1_rw_state(1), A2 => lbl1_rw_state(5), A3 => lbl1_rw_n_90, B1 => lbl1_rw_n_88, B2 => lbl1_rw_n_6, ZN => lbl1_rw_n_29);
  lbl1_rw_g2302 : IND3D1BWP7T port map(A1 => lbl1_n_1, B1 => go_to, B2 => FE_PHN53_lbl1_ready_rw, ZN => lbl1_rw_n_28);
  lbl1_rw_g2303 : AOI21D0BWP7T port map(A1 => lbl1_rw_n_86, A2 => lbl1_rw_state(1), B => lbl1_rw_n_85, ZN => lbl1_rw_n_27);
  lbl1_rw_g2304 : AOI21D0BWP7T port map(A1 => lbl1_rw_n_84, A2 => lbl1_rw_n_89, B => lbl1_rw_n_90, ZN => lbl1_rw_n_26);
  lbl1_rw_g2305 : CKXOR2D1BWP7T port map(A1 => write_memory(5), A2 => lbl1_cur_w(5), Z => lbl1_rw_n_25);
  lbl1_rw_g2306 : CKXOR2D1BWP7T port map(A1 => write_memory(7), A2 => lbl1_cur_w(7), Z => lbl1_rw_n_24);
  lbl1_rw_g2307 : CKXOR2D1BWP7T port map(A1 => write_memory(2), A2 => lbl1_cur_w(2), Z => lbl1_rw_n_23);
  lbl1_rw_g2308 : CKXOR2D1BWP7T port map(A1 => write_memory(1), A2 => lbl1_cur_w(1), Z => lbl1_rw_n_22);
  lbl1_rw_g2309 : CKXOR2D1BWP7T port map(A1 => write_memory(3), A2 => lbl1_cur_w(3), Z => lbl1_rw_n_21);
  lbl1_rw_g2310 : CKXOR2D1BWP7T port map(A1 => write_memory(0), A2 => lbl1_cur_w(0), Z => lbl1_rw_n_20);
  lbl1_rw_g2311 : CKXOR2D1BWP7T port map(A1 => address(6), A2 => y_address(1), Z => lbl1_rw_n_19);
  lbl1_rw_g2312 : CKXOR2D1BWP7T port map(A1 => address(1), A2 => x_address(1), Z => lbl1_rw_n_18);
  lbl1_rw_g2313 : CKXOR2D1BWP7T port map(A1 => address(7), A2 => y_address(2), Z => lbl1_rw_n_17);
  lbl1_rw_g2314 : XNR2D1BWP7T port map(A1 => address(9), A2 => y_address(4), ZN => lbl1_rw_n_16);
  lbl1_rw_g2315 : XNR2D1BWP7T port map(A1 => address(8), A2 => y_address(3), ZN => lbl1_rw_n_15);
  lbl1_rw_g2316 : CKXOR2D1BWP7T port map(A1 => address(2), A2 => x_address(2), Z => lbl1_rw_n_14);
  lbl1_rw_g2317 : CKXOR2D1BWP7T port map(A1 => address(5), A2 => y_address(0), Z => lbl1_rw_n_13);
  lbl1_rw_g2318 : XNR2D1BWP7T port map(A1 => address(0), A2 => x_address(0), ZN => lbl1_rw_n_12);
  lbl1_rw_g2319 : XNR2D1BWP7T port map(A1 => address(4), A2 => x_address(4), ZN => lbl1_rw_n_11);
  lbl1_rw_g2320 : XNR2D1BWP7T port map(A1 => address(3), A2 => x_address(3), ZN => lbl1_rw_n_10);
  lbl1_rw_g2321 : XNR2D1BWP7T port map(A1 => write_memory(6), A2 => lbl1_cur_w(6), ZN => lbl1_rw_n_9);
  lbl1_rw_g2322 : XNR2D1BWP7T port map(A1 => write_memory(4), A2 => lbl1_cur_w(4), ZN => lbl1_rw_n_8);
  lbl1_rw_g2323 : INVD0BWP7T port map(I => lbl1_rw_n_7, ZN => lbl1_rw_n_6);
  lbl1_rw_g2324 : CKND2D1BWP7T port map(A1 => lbl1_rw_state(0), A2 => lbl1_rw_state(4), ZN => lbl1_rw_n_7);
  lbl1_rw_g2325 : INVD0BWP7T port map(I => lbl1_rw_n_4, ZN => lbl1_rw_n_5);
  lbl1_rw_g2326 : OR2D1BWP7T port map(A1 => lbl1_rw_state(4), A2 => lbl1_rw_state(3), Z => lbl1_rw_n_3);
  lbl1_rw_g2327 : INR2XD0BWP7T port map(A1 => lbl1_rw_n_90, B1 => lbl1_rw_n_99, ZN => lbl1_rw_n_4);
  lbl1_rw_g2 : INR3D0BWP7T port map(A1 => lbl1_rw_n_43, B1 => lbl1_rw_n_7, B2 => FE_PHN83_lbl1_rw_state_2, ZN => lbl1_rw_n_0);
  lbl1_rw_state_reg_3 : DFD1BWP7T port map(CP => CTS_12, D => lbl1_rw_n_76, Q => lbl1_rw_state(3), QN => lbl1_rw_n_89);
  lbl1_rw_state_reg_5 : DFD1BWP7T port map(CP => CTS_12, D => FE_PHN69_lbl1_rw_n_60, Q => lbl1_rw_state(5), QN => lbl1_rw_n_87);
  lbl1_rw_state_reg_0 : DFD1BWP7T port map(CP => CTS_12, D => FE_PHN76_lbl1_rw_n_71, Q => lbl1_rw_state(0), QN => lbl1_rw_n_90);
  lbl1_rw_state_reg_1 : DFD1BWP7T port map(CP => CTS_12, D => lbl1_rw_n_74, Q => lbl1_rw_state(1), QN => lbl1_rw_n_88);
  lbl1_cey_g177 : OR2D1BWP7T port map(A1 => lbl1_cey_n_9, A2 => lbl1_cey_n_8, Z => lbl1_y_incr2);
  lbl1_cey_g178 : INR2D1BWP7T port map(A1 => lbl1_cey_state(1), B1 => lbl1_cey_state(0), ZN => lbl1_cey_n_8);
  lbl1_cey_g179 : INR2D1BWP7T port map(A1 => lbl1_cey_state(0), B1 => lbl1_cey_state(1), ZN => lbl1_cey_n_9);
  lbl1_cey_state_reg_0 : DFQD1BWP7T port map(CP => CTS_11, D => lbl1_cey_n_7, Q => lbl1_cey_state(0));
  lbl1_cey_g169 : NR2XD0BWP7T port map(A1 => FE_PHN73_lbl1_cey_n_6, A2 => FE_OFN3_rst, ZN => lbl1_cey_n_7);
  lbl1_cey_g171 : AOI21D0BWP7T port map(A1 => y_increment, A2 => lbl1_cey_n_4, B => lbl1_cey_n_8, ZN => lbl1_cey_n_6);
  lbl1_cey_g172 : NR2XD0BWP7T port map(A1 => lbl1_cey_n_3, A2 => FE_OFN3_rst, ZN => lbl1_cey_n_5);
  lbl1_cey_g173 : AOI21D0BWP7T port map(A1 => lbl1_n_1, A2 => lbl1_cey_n_2, B => lbl1_cey_n_9, ZN => lbl1_cey_n_4);
  lbl1_cey_g174 : AOI21D0BWP7T port map(A1 => y_increment, A2 => lbl1_cey_state(0), B => lbl1_y_incr2, ZN => FE_PHN71_lbl1_cey_n_3);
  lbl1_cey_state_reg_1 : DFD1BWP7T port map(CP => CTS_12, D => lbl1_cey_n_5, Q => lbl1_cey_state(1), QN => lbl1_cey_n_2);
  lbl1_cw_count_reg_7 : DFCNQD1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => w_increment_out, D => lbl1_cw_n_14, Q => lbl1_cur_w(7));
  lbl1_cw_g134 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_12, A2 => lbl1_cur_w(7), B1 => lbl1_cw_n_12, B2 => lbl1_cur_w(7), ZN => lbl1_cw_n_14);
  lbl1_cw_count_reg_6 : DFCNQD1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => w_increment_out, D => lbl1_cw_n_13, Q => lbl1_cur_w(6));
  lbl1_cw_g136 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_10, A2 => lbl1_cur_w(6), B1 => lbl1_cw_n_10, B2 => lbl1_cur_w(6), ZN => lbl1_cw_n_13);
  lbl1_cw_count_reg_5 : DFCNQD1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => w_increment_out, D => lbl1_cw_n_11, Q => lbl1_cur_w(5));
  lbl1_cw_g138 : IND2D0BWP7T port map(A1 => lbl1_cw_n_10, B1 => lbl1_cur_w(6), ZN => lbl1_cw_n_12);
  lbl1_cw_g139 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_8, A2 => lbl1_cur_w(5), B1 => lbl1_cw_n_8, B2 => lbl1_cur_w(5), ZN => lbl1_cw_n_11);
  lbl1_cw_count_reg_4 : DFCNQD1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => w_increment_out, D => lbl1_cw_n_9, Q => lbl1_cur_w(4));
  lbl1_cw_g141 : IND2D0BWP7T port map(A1 => lbl1_cw_n_8, B1 => lbl1_cur_w(5), ZN => lbl1_cw_n_10);
  lbl1_cw_g142 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_6, A2 => lbl1_cur_w(4), B1 => lbl1_cw_n_6, B2 => lbl1_cur_w(4), ZN => lbl1_cw_n_9);
  lbl1_cw_count_reg_3 : DFCNQD1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => w_increment_out, D => lbl1_cw_n_7, Q => lbl1_cur_w(3));
  lbl1_cw_g144 : IND2D0BWP7T port map(A1 => lbl1_cw_n_6, B1 => lbl1_cur_w(4), ZN => lbl1_cw_n_8);
  lbl1_cw_g145 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_4, A2 => lbl1_cur_w(3), B1 => lbl1_cw_n_4, B2 => lbl1_cur_w(3), ZN => lbl1_cw_n_7);
  lbl1_cw_count_reg_2 : DFCNQD1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => w_increment_out, D => lbl1_cw_n_5, Q => lbl1_cur_w(2));
  lbl1_cw_g147 : IND2D0BWP7T port map(A1 => lbl1_cw_n_4, B1 => lbl1_cur_w(3), ZN => lbl1_cw_n_6);
  lbl1_cw_g148 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_3, A2 => lbl1_cur_w(2), B1 => lbl1_cw_n_3, B2 => lbl1_cur_w(2), ZN => lbl1_cw_n_5);
  lbl1_cw_g150 : IND2D0BWP7T port map(A1 => lbl1_cw_n_3, B1 => lbl1_cur_w(2), ZN => lbl1_cw_n_4);
  lbl1_cw_g152 : ND2D0BWP7T port map(A1 => lbl1_cur_w(0), A2 => lbl1_cur_w(1), ZN => lbl1_cw_n_3);
  lbl1_cw_count_reg_0 : DFCND1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => w_increment_out, D => lbl1_cw_n_2, Q => lbl1_cur_w(0), QN => lbl1_cw_n_2);
  lbl1_cw_count_reg_1 : EDFCND1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => w_increment_out, D => lbl1_cw_n_0, E => lbl1_cur_w(0), Q => lbl1_cur_w(1), QN => lbl1_cw_n_0);
  lbl1_cx_count_reg_4 : DFCNQD1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => x_increment_out, D => lbl1_cx_n_8, Q => x_address(4));
  lbl1_cx_g82 : MOAI22D0BWP7T port map(A1 => lbl1_cx_n_6, A2 => x_address(4), B1 => lbl1_cx_n_6, B2 => x_address(4), ZN => lbl1_cx_n_8);
  lbl1_cx_count_reg_3 : DFCNQD1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => x_increment_out, D => lbl1_cx_n_7, Q => x_address(3));
  lbl1_cx_g84 : MOAI22D0BWP7T port map(A1 => lbl1_cx_n_4, A2 => x_address(3), B1 => lbl1_cx_n_4, B2 => x_address(3), ZN => lbl1_cx_n_7);
  lbl1_cx_count_reg_2 : DFCNQD1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => x_increment_out, D => lbl1_cx_n_5, Q => x_address(2));
  lbl1_cx_g86 : IND2D0BWP7T port map(A1 => lbl1_cx_n_4, B1 => x_address(3), ZN => lbl1_cx_n_6);
  lbl1_cx_g87 : MOAI22D0BWP7T port map(A1 => lbl1_cx_n_3, A2 => x_address(2), B1 => lbl1_cx_n_3, B2 => x_address(2), ZN => lbl1_cx_n_5);
  lbl1_cx_g89 : IND2D0BWP7T port map(A1 => lbl1_cx_n_3, B1 => x_address(2), ZN => lbl1_cx_n_4);
  lbl1_cx_g91 : ND2D0BWP7T port map(A1 => x_address(0), A2 => x_address(1), ZN => lbl1_cx_n_3);
  lbl1_cx_count_reg_1 : EDFCND1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => x_increment_out, D => lbl1_cx_n_2, E => x_address(0), Q => x_address(1), QN => lbl1_cx_n_2);
  lbl1_cx_count_reg_0 : DFCND1BWP7T port map(CDN => FE_DBTN3_memory_reset_out, CP => x_increment_out, D => lbl1_cx_n_0, Q => x_address(0), QN => lbl1_cx_n_0);
  lbl0_reg_n_layer_0_q_reg : EDFKCNQD1BWP7T port map(CN => FE_DBTN4_rst, CP => CTS_12, D => lbl0_n_474, E => lbl0_n_507, Q => lbl0_next_layer_0);

end routed;
