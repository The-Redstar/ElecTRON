library IEEE;
use IEEE.std_logic_1164.ALL;

entity countextend_tb is
end countextend_tb;

