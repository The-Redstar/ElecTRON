library IEEE;
use IEEE.std_logic_1164.ALL;

entity graphics_top_tb is
end graphics_top_tb;

