library IEEE;
use IEEE.std_logic_1164.ALL;

entity electron_tb is
end electron_tb;

