configuration test_data_gen_behaviour_cfg of test_data_gen is
   for behaviour
   end for;
end test_data_gen_behaviour_cfg;
