configuration electron_synthesised_cfg of electron is
   for synthesised
      for all: input_buffer use configuration work.input_buffer_behaviour_cfg;
      end for;
   end for;
end electron_synthesised_cfg;
