library IEEE;
use IEEE.std_logic_1164.ALL;

entity readwrite_tb is
end readwrite_tb;

