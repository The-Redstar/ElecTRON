configuration reg_3_behaviour_cfg of reg_3 is
   for behaviour
   end for;
end reg_3_behaviour_cfg;
