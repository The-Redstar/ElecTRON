library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of wall_decoder is
begin
end behaviour;

