library IEEE;
use IEEE.std_logic_1164.ALL;

entity counter8b_tb is
end counter8b_tb;

