library IEEE;
use IEEE.std_logic_1164.ALL;

entity sidebar_tb is
end sidebar_tb;

