configuration reg_1_behaviour_cfg of reg_1 is
   for behaviour
   end for;
end reg_1_behaviour_cfg;
