library IEEE;
use IEEE.std_logic_1164.ALL;

entity audio_top_tb is
end audio_top_tb;

