configuration graphics_top_tb_behaviour_cfg of graphics_top_tb is
   for behaviour
      for all: graphics_top use configuration work.graphics_top_behaviour_cfg;
      end for;
   end for;
end graphics_top_tb_behaviour_cfg;
