library IEEE;
use IEEE.std_logic_1164.ALL;

entity counter5b_tb is
end counter5b_tb;

