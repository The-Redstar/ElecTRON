library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity game_engine_tb is
end entity game_engine_tb;

architecture structural of game_engine_tb is

	component game_engine is
		port (clk                : in  std_logic;
        reset              : in  std_logic;
        input              : in  std_logic_vector(3 downto 0);
        busy               : in  std_logic;
        read_memory        : in  std_logic_vector(7 downto 0);
        memory_ready       : in  std_logic;
        state_vga          : out std_logic_vector(2 downto 0);
        write_enable       : out std_logic;
        write_memory       : out std_logic_vector(7 downto 0);
        address            : out std_logic_vector(9 downto 0);
        position_0_vga     : out std_logic_vector(10 downto 0);
        position_1_vga     : out std_logic_vector(10 downto 0);
        direction_0_vga    : out std_logic_vector(1 downto 0);
        direction_1_vga    : out std_logic_vector(1 downto 0);
        player_state_0_vga : out std_logic_vector(1 downto 0);
        player_state_1_vga : out std_logic_vector(1 downto 0);
		go_to	           : out std_logic;
		clear_memory       : out std_logic);
	end component game_engine;

	signal clk                : in  std_logic;
    signal reset              : in  std_logic;
    signal input              : in  std_logic_vector(3 downto 0);
    signal busy               : in  std_logic;
    signal read_memory        : in  std_logic_vector(7 downto 0);
    signal memory_ready       : in  std_logic;
    signal state_vga          : out std_logic_vector(2 downto 0);
    signal write_enable       : out std_logic;
    signal write_memory       : out std_logic_vector(7 downto 0);
    signal address            : out std_logic_vector(9 downto 0);
    signal position_0_vga     : out std_logic_vector(10 downto 0);
    signal position_1_vga     : out std_logic_vector(10 downto 0);
    signal direction_0_vga    : out std_logic_vector(1 downto 0);
    signal direction_1_vga    : out std_logic_vector(1 downto 0);
    signal player_state_0_vga : out std_logic_vector(1 downto 0);
    signal player_state_1_vga : out std_logic_vector(1 downto 0);
	signal go_to	          : out std_logic;
	signal clear_memory       : out std_logic;

begin

	lbl0: timebase port map	(clk               : clk,
							reset              : reset,
							input              : input,
							busy               : busy,
							read_memory        : read_memory,
							memory_ready       : memory_ready,
							state_vga          : state_vga,
							write_enable       : write_enable,
							write_memory       : write_memory,
							address            : address,
							position_0_vga     : position_0_vga,
							position_1_vga     : position_1_vga,
							direction_0_vga    : direction_0_vga,
							direction_1_vga    : direction_1_vga,
							player_state_0_vga : player_state_0_vga,
							player_state_1_vga : player_state_1_vga,
							go_to	           : go_to,
							clear_memory       : clear_memory
				);
					
end architecture structural;
