configuration reg_2_behaviour_cfg of reg_2 is
   for behaviour
   end for;
end reg_2_behaviour_cfg;
