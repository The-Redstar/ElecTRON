configuration input_buffer_behaviour_cfg of input_buffer is
   for behaviour
   end for;
end input_buffer_behaviour_cfg;
