configuration grid_top_behaviour_cfg of grid_top is
   for behaviour
   end for;
end grid_top_behaviour_cfg;
