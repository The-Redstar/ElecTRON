configuration sidebar_behaviour_cfg of sidebar is
   for behaviour
   end for;
end sidebar_behaviour_cfg;
