configuration graphics_top_behaviour_cfg of graphics_top is
   for behaviour
   end for;
end graphics_top_behaviour_cfg;
