
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture routed of electron is

  component DEL01BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL02BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL1BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD4BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD5BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD1BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD10BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component XNR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKXOR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component MOAI22D1BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component CKAN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKXOR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component DFD0BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component DFKSND1BWP7T
    port(CP, D, SN : in std_logic; Q, QN : out std_logic);
  end component;

  component DFKSND0BWP7T
    port(CP, D, SN : in std_logic; Q, QN : out std_logic);
  end component;

  component IINR4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD5BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AO222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component AO32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component IIND4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component DFXQD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component HA1D0BWP7T
    port(A, B : in std_logic; CO, S : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component INR4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component AOI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D1BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OA31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component OA32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component OR4XD1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component IND3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D2BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AO31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component IAO21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component XNR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component MUX2D1BWP7T
    port(I0, I1, S : in std_logic; Z : out std_logic);
  end component;

  component MAOI222D1BWP7T
    port(A, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OA221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component AN3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component OA222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component AO33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; Z : out std_logic);
  end component;

  component DFQD0BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component MUX2ND0BWP7T
    port(I0, I1, S : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D1BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component DFXD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q, QN : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component IOA21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AN4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component AN2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component FA1D0BWP7T
    port(A, B, CI : in std_logic; CO, S : out std_logic);
  end component;

  component OR3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component AN3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component OA22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component OA211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component OA33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; Z : out std_logic);
  end component;

  component OR3XD1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component MAOI22D1BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AN4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component AOI221D1BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component CKMUX2D1BWP7T
    port(I0, I1, S : in std_logic; Z : out std_logic);
  end component;

  component MUX2D0BWP7T
    port(I0, I1, S : in std_logic; Z : out std_logic);
  end component;

  component LNQD1BWP7T
    port(D, EN : in std_logic; Q : out std_logic);
  end component;

  component OR3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component OAI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component MAOI222D0BWP7T
    port(A, B, C : in std_logic; ZN : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AOI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component EDFKCNQD1BWP7T
    port(CN, CP, D, E : in std_logic; Q : out std_logic);
  end component;

  component OR3D4BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component CKAN2D8BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OR4D4BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component ND2D5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  signal FE_PHN349_lbl5_en1_new_period_17, FE_PHN348_lbl5_en1_new_period_1, FE_PHN347_lbl5_en1_new_period_3, FE_PHN346_lbl5_en1_n_10, FE_PHN345_lbl5_en1_new_period_5 : std_logic;
  signal FE_PHN344_lbl5_en1_n_301, FE_PHN343_lbl1_cm_n_8, FE_PHN342_lbl1_rw_n_84, FE_PHN341_lbl5_en0_new_period_6, FE_PHN340_lbl0_border_1 : std_logic;
  signal FE_PHN339_lbl1_cm_state_0, FE_PHN338_lbl5_en0_period_7, FE_PHN337_lbl5_en1_new_period_0, FE_PHN336_lbl2_v_count_7, FE_PHN335_lbl1_cur_w_1 : std_logic;
  signal FE_PHN334_lbl5_en1_new_period_4, FE_PHN333_lbl0_mem_com_state_2, FE_PHN332_lbl1_cur_w_3, FE_PHN331_lbl5_en1_new_period_5, FE_PHN330_lbl0_border_0 : std_logic;
  signal FE_PHN329_lbl5_en0_n_7, FE_PHN328_direction_in_2, FE_PHN327_lbl5_en1_n_3, FE_PHN326_lbl1_cur_w_5, FE_PHN325_lbl5_en1_count_6 : std_logic;
  signal FE_PHN324_y_address_0, FE_PHN323_lbl2_jumps_synced_7, FE_PHN322_lbl5_en1_new_period_17, FE_PHN321_lbl5_en1_new_period_1, FE_PHN320_lbl5_en1_n_10 : std_logic;
  signal FE_PHN319_lbl5_en1_new_period_3, FE_PHN318_lbl5_en0_new_period_5, FE_PHN317_lbl5_en1_new_period_14, FE_PHN316_lbl2_v_count_9, FE_PHN315_lbl0_busy_count_0 : std_logic;
  signal FE_PHN314_lbl0_mem_com_state_0, FE_PHN313_lbl5_en1_frozen_bits_1, FE_PHN312_lbl5_en1_new_period_8, FE_PHN311_lbl0_n_47, FE_PHN310_lbl1_cy_n_10 : std_logic;
  signal FE_PHN309_lbl0_n_539, FE_PHN308_lbl1_cm_n_23, FE_PHN307_lbl0_n_46, FE_PHN306_lbl5_en1_n_178, FE_PHN305_lbl1_cy_n_3 : std_logic;
  signal FE_PHN304_lbl1_cex_n_3, FE_PHN303_lbl1_cey_n_3, FE_PHN302_lbl1_cy_n_7, FE_PHN301_lbl1_cy_n_5, FE_PHN300_lbl1_cx_n_10 : std_logic;
  signal FE_PHN299_lbl1_cw_n_7, FE_PHN298_lbl1_cx_n_7, FE_PHN297_lbl1_cw_n_16, FE_PHN296_lbl1_cx_n_5, FE_PHN295_lbl5_expl_n_1 : std_logic;
  signal FE_PHN294_lbl0_n_34, FE_PHN293_lbl1_cm_n_24, FE_PHN292_lbl5_en0_n_46, FE_PHN291_lbl1_rw_n_68, FE_PHN290_lbl5_en1_n_300 : std_logic;
  signal FE_PHN289_lbl5_en1_n_179, FE_PHN288_lbl1_cw_n_3, FE_PHN287_lbl5_en1_n_183, FE_PHN286_lbl5_en0_n_296, FE_PHN285_lbl5_en0_n_157 : std_logic;
  signal FE_PHN284_lbl5_en0_n_156, FE_PHN283_lbl1_cx_n_3, FE_PHN282_lbl5_en0_n_161, FE_PHN281_lbl5_en0_n_298, FE_PHN280_lbl5_en1_n_302 : std_logic;
  signal FE_PHN279_lbl0_n_37, FE_PHN278_lbl5_en1_n_182, FE_PHN277_lbl1_cey_n_1, FE_PHN276_lbl0_n_43, FE_PHN275_lbl1_cex_n_1 : std_logic;
  signal FE_PHN274_lbl0_n_38, FE_PHN273_lbl5_en1_n_280, FE_PHN272_lbl0_n_42, FE_PHN271_lbl5_en0_n_276, FE_PHN270_lbl5_en0_n_155 : std_logic;
  signal FE_PHN269_lbl0_n_45, FE_PHN268_lbl0_n_44, FE_PHN267_lbl5_en0_n_158, FE_PHN266_lbl0_mem_com_state_0, FE_PHN265_lbl5_en0_new_period_6 : std_logic;
  signal FE_PHN264_lbl5_en0_period_18, FE_PHN263_lbl5_en0_period_16, FE_PHN262_lbl0_mem_com_state_3, FE_PHN261_lbl5_en0_period_17, FE_PHN260_lbl5_en1_period_17 : std_logic;
  signal FE_PHN259_lbl5_en1_period_16, FE_PHN258_lbl0_busy_count_0, FE_PHN257_x_address_3, FE_PHN256_lbl0_mem_com_state_1, FE_PHN255_direction_0_1 : std_logic;
  signal FE_PHN254_lbl5_en0_count_16, FE_PHN253_direction_between_3, FE_PHN252_lbl5_en1_new_period_1, FE_PHN251_lbl5_en0_count_17, FE_PHN250_lbl5_en1_new_period_5 : std_logic;
  signal FE_PHN249_lbl5_en0_new_period_5, FE_PHN248_lbl5_en1_new_period_3, FE_PHN247_y_address_3, FE_PHN246_lbl5_en0_new_period_2, FE_PHN245_lbl5_en1_n_10 : std_logic;
  signal FE_PHN244_lbl5_en1_new_period_2, FE_PHN243_lbl5_en0_new_period_14, FE_PHN242_lbl5_en0_new_period_4, FE_PHN241_direction_between_2, FE_PHN240_direction_between_0 : std_logic;
  signal FE_PHN239_lbl5_en1_new_period_7, FE_PHN238_lbl2_v_count_9, FE_PHN237_lbl5_en0_new_period_8, FE_PHN236_lbl5_en0_new_period_13, FE_PHN235_read_memory_in_4 : std_logic;
  signal FE_PHN234_lbl5_en0_new_period_10, FE_PHN233_lbl5_en0_new_period_11, FE_PHN232_lbl5_en0_n_7, FE_PHN231_read_memory_in_5, FE_PHN230_lbl5_en0_new_period_9 : std_logic;
  signal FE_PHN229_lbl2_n_21, FE_PHN228_lbl5_en1_new_period_13, FE_PHN227_lbl5_en1_n_4, FE_PHN226_lbl5_en1_n_2, FE_PHN225_lbl5_en1_new_period_4 : std_logic;
  signal FE_PHN224_lbl5_en1_n_3, FE_PHN223_lbl5_en1_n_8, FE_PHN222_lbl5_en1_n_9, FE_PHN221_lbl5_en1_new_period_14, FE_PHN220_lbl5_en0_new_period_7 : std_logic;
  signal FE_PHN219_lbl5_en0_new_period_0, FE_PHN218_direction_between_1, FE_PHN217_read_memory_in_0, FE_PHN216_lbl5_en1_new_period_8, FE_PHN215_lbl5_en1_new_period_9 : std_logic;
  signal FE_PHN214_lbl1_cur_w_1, FE_PHN213_lbl5_en1_new_period_16, FE_PHN212_lbl1_cur_w_2, FE_PHN211_lbl5_en1_new_period_0, FE_PHN210_lbl0_n_65 : std_logic;
  signal FE_PHN209_lbl5_en1_n_6, FE_PHN208_lbl1_cur_w_3, FE_PHN207_lbl0_n_81, FE_PHN206_lbl5_en1_new_period_11, FE_PHN205_read_memory_in_1 : std_logic;
  signal FE_PHN204_lbl5_en1_n_7, FE_PHN203_lbl5_en1_new_period_15, FE_PHN202_lbl5_en0_new_period_15, FE_PHN201_read_memory_in_2, FE_PHN200_lbl1_cur_w_0 : std_logic;
  signal FE_PHN199_lbl5_en0_frozen_boost, FE_PHN198_read_memory_in_6, FE_PHN197_lbl1_cur_w_4, FE_PHN196_lbl0_next_direction_0_1, FE_PHN195_lbl5_en1_n_290 : std_logic;
  signal FE_PHN194_lbl2_v_count_7, FE_PHN193_read_memory_in_7, FE_PHN192_lbl5_en0_new_period_16, FE_PHN191_lbl1_cur_w_6, FE_PHN190_lbl5_en1_n_285 : std_logic;
  signal FE_PHN189_lbl5_en1_n_292, FE_PHN188_lbl5_en0_n_281, FE_PHN187_lbl1_cur_w_5, FE_PHN186_lbl1_rw_n_0, FE_PHN185_lbl5_en1_count_17 : std_logic;
  signal FE_PHN184_lbl5_en0_n_285, FE_PHN183_lbl5_en1_n_288, FE_PHN182_lbl0_counter_busy_counter_state_0, FE_PHN181_lbl5_en0_n_283, FE_PHN180_lbl5_en0_n_289 : std_logic;
  signal FE_PHN179_lbl5_en1_n_287, FE_PHN178_lbl5_en1_n_289, FE_PHN177_lbl5_en0_n_282, FE_PHN176_lbl5_en0_n_290, FE_PHN175_lbl5_en0_n_291 : std_logic;
  signal FE_PHN174_lbl1_cm_n_52, FE_PHN173_lbl5_en1_n_293, FE_PHN172_lbl5_en0_n_293, FE_PHN171_direction_0_0, FE_PHN170_lbl5_en1_n_295 : std_logic;
  signal FE_PHN169_lbl5_en0_n_288, FE_PHN168_lbl5_en0_n_287, FE_PHN167_lbl0_n_63, FE_PHN166_lbl5_en0_n_286, FE_PHN165_lbl5_en0_n_284 : std_logic;
  signal FE_PHN164_lbl0_counter_busy_counter_state_1, FE_PHN163_lbl0_border_0, FE_PHN162_lbl5_en1_n_298, FE_PHN161_lbl5_en1_n_294, FE_PHN160_lbl5_en0_n_292 : std_logic;
  signal FE_PHN159_lbl5_en1_n_291, FE_PHN158_lbl5_en0_n_294, FE_PHN157_lbl1_cex_n_4, FE_PHN156_lbl1_cm_n_22, FE_PHN155_lbl0_border_1 : std_logic;
  signal FE_PHN154_lbl1_cey_n_4, FE_PHN153_read_memory_in_3, FE_PHN152_lbl1_rw_n_27, FE_PHN151_direction_in_2, FE_PHN150_lbl2_v_count_8 : std_logic;
  signal FE_PHN149_lbl1_rw_n_58, FE_PHN148_lbl5_en1_n_296, FE_PHN147_lbl5_en1_period_4, FE_PHN146_lbl5_en1_n_5, FE_PHN145_lbl5_en0_period_7 : std_logic;
  signal FE_PHN144_lbl5_en0_period_13, FE_PHN143_lbl2_jumps_synced_7, FE_PHN142_boost_audio_1, FE_PHN141_lbl5_en0_n_295, FE_PHN140_lbl5_en1_frozen_boost : std_logic;
  signal FE_PHN139_lbl5_en1_n_299, FE_PHN138_lbl2_v_count_6, FE_PHN137_lbl5_en1_count_16, FE_PHN136_lbl5_en1_new_period_17, FE_PHN135_lbl5_en1_n_297 : std_logic;
  signal FE_PHN134_direction_in_0, FE_PHN133_lbl2_data_synced_2, FE_PHN132_lbl5_en0_period_10, FE_PHN131_lbl5_en1_frozen_bits_0, FE_PHN130_lbl5_en1_n_286 : std_logic;
  signal FE_PHN129_lbl2_data_synced_1, FE_PHN128_direction_1_1, FE_PHN127_direction_in_1, FE_PHN126_direction_1_0, FE_PHN125_lbl5_en1_frozen_bits_1 : std_logic;
  signal FE_PHN124_lbl5_en0_period_5, FE_PHN123_lbl5_en1_period_6, FE_PHN122_lbl2_data_synced_5, FE_PHN121_lbl5_en0_frozen_bits_2, FE_PHN120_lbl2_data_synced_6 : std_logic;
  signal FE_PHN119_lbl5_en1_period_5, FE_PHN118_lbl5_en0_n_6, FE_PHN117_lbl5_en1_n_13, FE_PHN116_lbl2_data_synced_0, FE_PHN115_lbl5_en0_period_9 : std_logic;
  signal FE_PHN114_lbl5_en1_period_9, FE_PHN113_lbl5_en1_period_7, FE_PHN112_lbl5_en1_period_12, FE_PHN111_lbl5_en0_n_8, FE_PHN110_lbl5_en0_period_3 : std_logic;
  signal FE_PHN109_lbl2_data_synced_4, FE_PHN108_lbl5_en0_frozen_bits_3, FE_PHN107_lbl5_en0_period_14, FE_PHN106_lbl5_en1_period_10, FE_PHN105_lbl5_en0_period_12 : std_logic;
  signal FE_PHN104_boost_audio_0, FE_PHN103_direction_in_3, FE_PHN102_lbl5_en1_period_11, FE_PHN101_lbl2_data_synced_3, FE_PHN100_lbl5_en0_n_5 : std_logic;
  signal FE_PHN99_lbl5_en1_period_1, FE_PHN98_lbl5_en0_period_2, FE_PHN97_lbl5_en0_period_8, FE_PHN96_lbl5_en1_frozen_bits_3, FE_PHN95_lbl5_en1_period_13 : std_logic;
  signal FE_PHN94_lbl2_borders_synced_1, FE_PHN93_lbl2_borders_synced_5, FE_PHN92_lbl5_en0_period_6, FE_PHN91_lbl5_en0_period_15, FE_PHN90_lbl5_en1_period_14 : std_logic;
  signal FE_PHN89_lbl5_en1_period_8, FE_PHN88_lbl5_en0_period_0, FE_PHN87_lbl5_en1_period_18, FE_PHN86_lbl5_en1_period_0, FE_PHN85_lbl2_borders_synced_6 : std_logic;
  signal FE_PHN84_lbl5_en1_period_15, FE_PHN83_lbl2_borders_synced_2, FE_PHN82_lbl2_borders_synced_7, FE_PHN81_lbl5_en1_frozen_bits_2, FE_PHN80_lbl5_en0_period_4 : std_logic;
  signal FE_PHN79_lbl2_data_synced_7, FE_PHN78_lbl2_jumps_synced_5, FE_PHN77_lbl2_jumps_synced_3, FE_PHN76_lbl2_jumps_synced_6, FE_PHN75_lbl2_jumps_synced_0 : std_logic;
  signal FE_PHN74_lbl2_borders_synced_4, FE_PHN73_lbl2_borders_synced_3, FE_PHN72_lbl5_en0_period_11, FE_PHN71_lbl2_jumps_synced_1, FE_PHN70_lbl5_en1_period_2 : std_logic;
  signal FE_PHN69_lbl2_jumps_synced_4, FE_PHN68_lbl2_borders_synced_0, FE_PHN67_lbl2_jumps_synced_2, FE_PHN66_lbl5_en1_period_3, FE_PHN65_start_in : std_logic;
  signal FE_PHN64_lbl5_en0_new_period_17, FE_PHN63_lbl5_en0_period_1, FE_PHN62_lbl5_en0_n_12, FE_PHN61_lbl0_booster_sync, FE_PHN60_lbl5_expl_shifter_15 : std_logic;
  signal FE_PHN59_lbl5_expl_shifter_21, FE_PHN58_lbl5_expl_shifter_6, FE_PHN57_lbl5_en0_frozen_bits_0, FE_PHN56_lbl5_en0_n_16, FE_PHN55_lbl3_temp1_1 : std_logic;
  signal FE_PHN54_lbl5_en0_n_11, FE_PHN53_lbl5_en0_frozen_bits_1, FE_PHN52_lbl5_en0_n_14, FE_PHN51_lbl5_en0_n_9, FE_PHN50_lbl3_temp2 : std_logic;
  signal FE_PHN49_lbl5_expl_shifter_20, FE_PHN48_lbl3_temp1_0, FE_PHN47_lbl5_expl_shifter_4, FE_PHN46_lbl5_expl_shifter_22, FE_PHN45_lbl5_expl_shifter_17 : std_logic;
  signal FE_PHN44_lbl5_expl_shifter_16, FE_PHN43_lbl5_expl_shifter_7, FE_PHN42_lbl5_expl_shifter_5, FE_PHN41_lbl5_expl_shifter_13, FE_PHN40_lbl5_expl_shifter_11 : std_logic;
  signal FE_PHN39_lbl5_expl_shifter_14, FE_PHN38_lbl5_expl_shifter_10, FE_PHN37_lbl5_expl_shifter_12, FE_PHN36_lbl5_expl_shifter_9, FE_PHN35_lbl5_expl_shifter_8 : std_logic;
  signal FE_PHN34_lbl5_expl_shifter_18, FE_PHN33_lbl5_expl_shifter_19, FE_PHN32_lbl3_temp1_3, FE_PHN31_lbl5_en1_new_period_18, FE_PHN30_lbl5_en0_new_period_18 : std_logic;
  signal FE_PHN29_lbl3_temp1_2, FE_PHN28_lbl5_bits_3, FE_PHN27_lbl5_bits_2, FE_PHN26_lbl5_bits_0, FE_PHN25_lbl5_bits_1 : std_logic;
  signal FE_OFN5_FE_DBTN24_rst, FE_OFN4_memory_enable_out, FE_OFN1_rst, FE_OFN0_lbl2_n_2, CTS_22 : std_logic;
  signal CTS_21, CTS_20, CTS_19, CTS_18, FE_DBTN24_rst : std_logic;
  signal FE_DBTN23_memory_reset_out, FE_DBTN22_position_1_10, FE_DBTN21_lbl2_h_count_3, FE_DBTN20_lbl2_h_count_2, FE_DBTN19_lbl2_h_count_1 : std_logic;
  signal FE_DBTN18_lbl2_v_count_2, FE_DBTN17_lbl5_en0_n_301, FE_DBTN16_lbl5_en0_n_304, FE_DBTN15_lbl5_en0_n_306, FE_DBTN14_lbl5_en0_n_305 : std_logic;
  signal FE_DBTN13_lbl5_en0_n_309, FE_DBTN12_lbl5_en0_n_303, FE_DBTN11_lbl5_en0_n_308, FE_DBTN10_lbl5_en0_n_311, FE_DBTN9_lbl5_en0_n_302 : std_logic;
  signal FE_DBTN8_lbl5_en1_n_305, FE_DBTN7_lbl5_en1_n_308, FE_DBTN6_lbl5_en1_n_310, FE_DBTN5_lbl5_en1_n_309, FE_DBTN4_lbl5_en1_n_313 : std_logic;
  signal FE_DBTN3_lbl5_en1_n_307, FE_DBTN2_lbl5_en1_n_312, FE_DBTN1_lbl5_en1_n_315, FE_DBTN0_lbl5_en1_n_306 : std_logic;
  signal position_1 : std_logic_vector(10 downto 0);
  signal position_0 : std_logic_vector(10 downto 0);
  signal lbl2_y_vec : std_logic_vector(4 downto 0);
  signal lbl2_central_x_vec : std_logic_vector(9 downto 0);
  signal lbl2_h_count : std_logic_vector(9 downto 0);
  signal lbl2_dx : std_logic_vector(3 downto 0);
  signal lbl2_v_count : std_logic_vector(9 downto 0);
  signal lbl2_dy_vec : std_logic_vector(3 downto 0);
  signal game_state : std_logic_vector(2 downto 0);
  signal lbl2_homescreen_color : std_logic_vector(3 downto 0);
  signal lbl2_pixelator_color : std_logic_vector(3 downto 0);
  signal lbl2_sidebar_color : std_logic_vector(3 downto 0);
  signal direction_between : std_logic_vector(3 downto 0);
  signal player_state_0 : std_logic_vector(1 downto 0);
  signal player_state_1 : std_logic_vector(1 downto 0);
  signal lbl2_borders_synced : std_logic_vector(7 downto 0);
  signal borders : std_logic_vector(7 downto 0);
  signal lbl2_data_synced : std_logic_vector(7 downto 0);
  signal lbl2_jumps_synced : std_logic_vector(7 downto 0);
  signal ramps : std_logic_vector(7 downto 0);
  signal lbl3_temp1 : std_logic_vector(3 downto 0);
  signal lbl2_walls : std_logic_vector(7 downto 0);
  signal x_address : std_logic_vector(4 downto 0);
  signal start_position_0 : std_logic_vector(10 downto 0);
  signal y_address : std_logic_vector(4 downto 0);
  signal map_selected : std_logic_vector(1 downto 0);
  signal start_position_1 : std_logic_vector(10 downto 0);
  signal lbl5_expl_shifter : std_logic_vector(23 downto 0);
  signal lbl5_bits : std_logic_vector(3 downto 0);
  signal lbl5_en0_period : std_logic_vector(18 downto 0);
  signal direction_0 : std_logic_vector(1 downto 0);
  signal lbl5_en0_prev_dir : std_logic_vector(1 downto 0);
  signal lbl5_en0_frozen_bits : std_logic_vector(3 downto 0);
  signal lbl5_en0_count : std_logic_vector(18 downto 0);
  signal lbl5_en0_new_period : std_logic_vector(18 downto 0);
  signal lbl5_en1_period : std_logic_vector(18 downto 0);
  signal direction_1 : std_logic_vector(1 downto 0);
  signal lbl5_en1_prev_dir : std_logic_vector(1 downto 0);
  signal lbl5_en1_frozen_bits : std_logic_vector(3 downto 0);
  signal lbl5_en1_count : std_logic_vector(18 downto 0);
  signal lbl5_en1_new_period : std_logic_vector(18 downto 0);
  signal lbl0_new_state : std_logic_vector(4 downto 0);
  signal lbl0_d_position_1 : std_logic_vector(9 downto 0);
  signal address : std_logic_vector(9 downto 0);
  signal lbl0_next_direction_0 : std_logic_vector(1 downto 0);
  signal lbl0_next_direction_1 : std_logic_vector(1 downto 0);
  signal lbl0_d_position_0 : std_logic_vector(9 downto 0);
  signal lbl0_d_read_data_reg : std_logic_vector(7 downto 0);
  signal lbl0_busy_count : std_logic_vector(6 downto 0);
  signal lbl0_state : std_logic_vector(4 downto 0);
  signal write_memory : std_logic_vector(7 downto 0);
  signal lbl0_read_data_reg : std_logic_vector(7 downto 0);
  signal lbl0_mem_com_state : std_logic_vector(3 downto 0);
  signal lbl0_d_next_direction_1 : std_logic_vector(1 downto 0);
  signal lbl0_d_next_direction_0 : std_logic_vector(1 downto 0);
  signal lbl0_d_speed_select : std_logic_vector(1 downto 0);
  signal lbl0_d_map_select : std_logic_vector(1 downto 0);
  signal lbl0_d_direction_0 : std_logic_vector(1 downto 0);
  signal lbl0_d_direction_1 : std_logic_vector(1 downto 0);
  signal lbl0_counter_busy_counter_state : std_logic_vector(1 downto 0);
  signal lbl1_cm_state : std_logic_vector(4 downto 0);
  signal lbl1_cex_state : std_logic_vector(1 downto 0);
  signal lbl1_rw_state : std_logic_vector(5 downto 0);
  signal lbl1_cur_w : std_logic_vector(7 downto 0);
  signal lbl1_cey_state : std_logic_vector(1 downto 0);
  signal UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2, UNCONNECTED3 : std_logic;
  signal UNCONNECTED4, UNCONNECTED5, UNCONNECTED6, UNCONNECTED7, UNCONNECTED8 : std_logic;
  signal UNCONNECTED9, boost_audio_0, boost_audio_1, busy, clear_memory : std_logic;
  signal go_to, lbl0_booster_sync, lbl0_border_0, lbl0_border_1, lbl0_d_booster_sync : std_logic;
  signal lbl0_d_layer_0, lbl0_d_layer_1, lbl0_d_move_0, lbl0_d_move_1, lbl0_e_position_0 : std_logic;
  signal lbl0_e_position_1, lbl0_mem_com_n_166, lbl0_mem_com_n_175, lbl0_move_0, lbl0_move_1 : std_logic;
  signal lbl0_n_0, lbl0_n_1, lbl0_n_2, lbl0_n_4, lbl0_n_5 : std_logic;
  signal lbl0_n_6, lbl0_n_7, lbl0_n_9, lbl0_n_10, lbl0_n_11 : std_logic;
  signal lbl0_n_12, lbl0_n_13, lbl0_n_14, lbl0_n_15, lbl0_n_16 : std_logic;
  signal lbl0_n_17, lbl0_n_18, lbl0_n_19, lbl0_n_20, lbl0_n_21 : std_logic;
  signal lbl0_n_22, lbl0_n_23, lbl0_n_24, lbl0_n_25, lbl0_n_27 : std_logic;
  signal lbl0_n_28, lbl0_n_30, lbl0_n_31, lbl0_n_32, lbl0_n_33 : std_logic;
  signal lbl0_n_34, lbl0_n_35, lbl0_n_36, lbl0_n_37, lbl0_n_38 : std_logic;
  signal lbl0_n_40, lbl0_n_41, lbl0_n_42, lbl0_n_43, lbl0_n_44 : std_logic;
  signal lbl0_n_45, lbl0_n_46, lbl0_n_47, lbl0_n_48, lbl0_n_49 : std_logic;
  signal lbl0_n_50, lbl0_n_51, lbl0_n_52, lbl0_n_53, lbl0_n_54 : std_logic;
  signal lbl0_n_55, lbl0_n_56, lbl0_n_58, lbl0_n_59, lbl0_n_60 : std_logic;
  signal lbl0_n_61, lbl0_n_62, lbl0_n_63, lbl0_n_64, lbl0_n_65 : std_logic;
  signal lbl0_n_66, lbl0_n_67, lbl0_n_68, lbl0_n_71, lbl0_n_72 : std_logic;
  signal lbl0_n_73, lbl0_n_74, lbl0_n_75, lbl0_n_76, lbl0_n_78 : std_logic;
  signal lbl0_n_79, lbl0_n_80, lbl0_n_81, lbl0_n_82, lbl0_n_83 : std_logic;
  signal lbl0_n_84, lbl0_n_85, lbl0_n_86, lbl0_n_87, lbl0_n_88 : std_logic;
  signal lbl0_n_89, lbl0_n_90, lbl0_n_91, lbl0_n_92, lbl0_n_93 : std_logic;
  signal lbl0_n_94, lbl0_n_95, lbl0_n_96, lbl0_n_97, lbl0_n_98 : std_logic;
  signal lbl0_n_99, lbl0_n_100, lbl0_n_101, lbl0_n_102, lbl0_n_103 : std_logic;
  signal lbl0_n_104, lbl0_n_105, lbl0_n_106, lbl0_n_107, lbl0_n_108 : std_logic;
  signal lbl0_n_109, lbl0_n_110, lbl0_n_111, lbl0_n_112, lbl0_n_113 : std_logic;
  signal lbl0_n_114, lbl0_n_115, lbl0_n_116, lbl0_n_117, lbl0_n_118 : std_logic;
  signal lbl0_n_119, lbl0_n_120, lbl0_n_121, lbl0_n_122, lbl0_n_123 : std_logic;
  signal lbl0_n_124, lbl0_n_125, lbl0_n_126, lbl0_n_127, lbl0_n_128 : std_logic;
  signal lbl0_n_129, lbl0_n_130, lbl0_n_131, lbl0_n_132, lbl0_n_133 : std_logic;
  signal lbl0_n_134, lbl0_n_135, lbl0_n_136, lbl0_n_137, lbl0_n_138 : std_logic;
  signal lbl0_n_139, lbl0_n_140, lbl0_n_141, lbl0_n_142, lbl0_n_143 : std_logic;
  signal lbl0_n_144, lbl0_n_145, lbl0_n_146, lbl0_n_147, lbl0_n_148 : std_logic;
  signal lbl0_n_149, lbl0_n_150, lbl0_n_151, lbl0_n_152, lbl0_n_153 : std_logic;
  signal lbl0_n_154, lbl0_n_155, lbl0_n_156, lbl0_n_157, lbl0_n_158 : std_logic;
  signal lbl0_n_159, lbl0_n_160, lbl0_n_161, lbl0_n_162, lbl0_n_163 : std_logic;
  signal lbl0_n_164, lbl0_n_165, lbl0_n_166, lbl0_n_167, lbl0_n_168 : std_logic;
  signal lbl0_n_169, lbl0_n_170, lbl0_n_171, lbl0_n_172, lbl0_n_173 : std_logic;
  signal lbl0_n_174, lbl0_n_175, lbl0_n_176, lbl0_n_177, lbl0_n_178 : std_logic;
  signal lbl0_n_179, lbl0_n_180, lbl0_n_181, lbl0_n_182, lbl0_n_183 : std_logic;
  signal lbl0_n_184, lbl0_n_185, lbl0_n_186, lbl0_n_187, lbl0_n_188 : std_logic;
  signal lbl0_n_189, lbl0_n_190, lbl0_n_191, lbl0_n_192, lbl0_n_193 : std_logic;
  signal lbl0_n_194, lbl0_n_195, lbl0_n_196, lbl0_n_197, lbl0_n_198 : std_logic;
  signal lbl0_n_199, lbl0_n_200, lbl0_n_201, lbl0_n_202, lbl0_n_203 : std_logic;
  signal lbl0_n_204, lbl0_n_205, lbl0_n_206, lbl0_n_207, lbl0_n_208 : std_logic;
  signal lbl0_n_209, lbl0_n_210, lbl0_n_211, lbl0_n_212, lbl0_n_213 : std_logic;
  signal lbl0_n_214, lbl0_n_215, lbl0_n_216, lbl0_n_217, lbl0_n_218 : std_logic;
  signal lbl0_n_219, lbl0_n_220, lbl0_n_221, lbl0_n_222, lbl0_n_223 : std_logic;
  signal lbl0_n_224, lbl0_n_225, lbl0_n_226, lbl0_n_227, lbl0_n_228 : std_logic;
  signal lbl0_n_229, lbl0_n_230, lbl0_n_231, lbl0_n_232, lbl0_n_233 : std_logic;
  signal lbl0_n_234, lbl0_n_235, lbl0_n_236, lbl0_n_237, lbl0_n_238 : std_logic;
  signal lbl0_n_239, lbl0_n_240, lbl0_n_241, lbl0_n_242, lbl0_n_243 : std_logic;
  signal lbl0_n_244, lbl0_n_245, lbl0_n_246, lbl0_n_247, lbl0_n_248 : std_logic;
  signal lbl0_n_249, lbl0_n_250, lbl0_n_251, lbl0_n_252, lbl0_n_253 : std_logic;
  signal lbl0_n_254, lbl0_n_255, lbl0_n_256, lbl0_n_257, lbl0_n_258 : std_logic;
  signal lbl0_n_259, lbl0_n_260, lbl0_n_261, lbl0_n_262, lbl0_n_263 : std_logic;
  signal lbl0_n_264, lbl0_n_265, lbl0_n_266, lbl0_n_267, lbl0_n_268 : std_logic;
  signal lbl0_n_269, lbl0_n_270, lbl0_n_271, lbl0_n_272, lbl0_n_273 : std_logic;
  signal lbl0_n_274, lbl0_n_275, lbl0_n_276, lbl0_n_277, lbl0_n_278 : std_logic;
  signal lbl0_n_279, lbl0_n_280, lbl0_n_281, lbl0_n_282, lbl0_n_283 : std_logic;
  signal lbl0_n_284, lbl0_n_285, lbl0_n_286, lbl0_n_287, lbl0_n_288 : std_logic;
  signal lbl0_n_289, lbl0_n_290, lbl0_n_291, lbl0_n_292, lbl0_n_293 : std_logic;
  signal lbl0_n_294, lbl0_n_295, lbl0_n_296, lbl0_n_297, lbl0_n_298 : std_logic;
  signal lbl0_n_299, lbl0_n_300, lbl0_n_301, lbl0_n_302, lbl0_n_303 : std_logic;
  signal lbl0_n_304, lbl0_n_305, lbl0_n_306, lbl0_n_307, lbl0_n_308 : std_logic;
  signal lbl0_n_309, lbl0_n_310, lbl0_n_311, lbl0_n_312, lbl0_n_313 : std_logic;
  signal lbl0_n_314, lbl0_n_315, lbl0_n_316, lbl0_n_317, lbl0_n_318 : std_logic;
  signal lbl0_n_319, lbl0_n_320, lbl0_n_321, lbl0_n_322, lbl0_n_323 : std_logic;
  signal lbl0_n_324, lbl0_n_325, lbl0_n_326, lbl0_n_327, lbl0_n_328 : std_logic;
  signal lbl0_n_329, lbl0_n_330, lbl0_n_331, lbl0_n_332, lbl0_n_333 : std_logic;
  signal lbl0_n_334, lbl0_n_335, lbl0_n_336, lbl0_n_337, lbl0_n_338 : std_logic;
  signal lbl0_n_339, lbl0_n_340, lbl0_n_341, lbl0_n_342, lbl0_n_343 : std_logic;
  signal lbl0_n_345, lbl0_n_346, lbl0_n_347, lbl0_n_348, lbl0_n_349 : std_logic;
  signal lbl0_n_350, lbl0_n_351, lbl0_n_352, lbl0_n_353, lbl0_n_354 : std_logic;
  signal lbl0_n_355, lbl0_n_356, lbl0_n_357, lbl0_n_358, lbl0_n_359 : std_logic;
  signal lbl0_n_360, lbl0_n_361, lbl0_n_362, lbl0_n_363, lbl0_n_364 : std_logic;
  signal lbl0_n_365, lbl0_n_366, lbl0_n_367, lbl0_n_368, lbl0_n_369 : std_logic;
  signal lbl0_n_370, lbl0_n_371, lbl0_n_372, lbl0_n_373, lbl0_n_374 : std_logic;
  signal lbl0_n_375, lbl0_n_376, lbl0_n_377, lbl0_n_378, lbl0_n_379 : std_logic;
  signal lbl0_n_380, lbl0_n_381, lbl0_n_382, lbl0_n_383, lbl0_n_384 : std_logic;
  signal lbl0_n_385, lbl0_n_386, lbl0_n_387, lbl0_n_388, lbl0_n_389 : std_logic;
  signal lbl0_n_390, lbl0_n_391, lbl0_n_392, lbl0_n_393, lbl0_n_394 : std_logic;
  signal lbl0_n_395, lbl0_n_396, lbl0_n_397, lbl0_n_398, lbl0_n_399 : std_logic;
  signal lbl0_n_400, lbl0_n_401, lbl0_n_402, lbl0_n_403, lbl0_n_404 : std_logic;
  signal lbl0_n_405, lbl0_n_406, lbl0_n_407, lbl0_n_408, lbl0_n_409 : std_logic;
  signal lbl0_n_410, lbl0_n_411, lbl0_n_412, lbl0_n_413, lbl0_n_414 : std_logic;
  signal lbl0_n_415, lbl0_n_416, lbl0_n_417, lbl0_n_418, lbl0_n_419 : std_logic;
  signal lbl0_n_420, lbl0_n_421, lbl0_n_422, lbl0_n_423, lbl0_n_424 : std_logic;
  signal lbl0_n_425, lbl0_n_426, lbl0_n_427, lbl0_n_428, lbl0_n_429 : std_logic;
  signal lbl0_n_430, lbl0_n_431, lbl0_n_432, lbl0_n_433, lbl0_n_434 : std_logic;
  signal lbl0_n_436, lbl0_n_437, lbl0_n_438, lbl0_n_439, lbl0_n_440 : std_logic;
  signal lbl0_n_441, lbl0_n_442, lbl0_n_443, lbl0_n_444, lbl0_n_445 : std_logic;
  signal lbl0_n_446, lbl0_n_447, lbl0_n_448, lbl0_n_449, lbl0_n_450 : std_logic;
  signal lbl0_n_451, lbl0_n_452, lbl0_n_453, lbl0_n_454, lbl0_n_455 : std_logic;
  signal lbl0_n_456, lbl0_n_457, lbl0_n_461, lbl0_n_497, lbl0_n_498 : std_logic;
  signal lbl0_n_499, lbl0_n_500, lbl0_n_502, lbl0_n_503, lbl0_n_530 : std_logic;
  signal lbl0_n_531, lbl0_n_532, lbl0_n_533, lbl0_n_535, lbl0_n_536 : std_logic;
  signal lbl0_n_539, lbl0_n_541, lbl0_n_542, lbl0_next_layer_0, lbl0_next_layer_1 : std_logic;
  signal lbl1_cex_n_0, lbl1_cex_n_1, lbl1_cex_n_2, lbl1_cex_n_3, lbl1_cex_n_4 : std_logic;
  signal lbl1_cex_n_5, lbl1_cey_n_0, lbl1_cey_n_1, lbl1_cey_n_2, lbl1_cey_n_3 : std_logic;
  signal lbl1_cey_n_4, lbl1_cey_n_5, lbl1_clr_rst, lbl1_cm_n_0, lbl1_cm_n_1 : std_logic;
  signal lbl1_cm_n_2, lbl1_cm_n_3, lbl1_cm_n_4, lbl1_cm_n_5, lbl1_cm_n_6 : std_logic;
  signal lbl1_cm_n_7, lbl1_cm_n_8, lbl1_cm_n_9, lbl1_cm_n_11, lbl1_cm_n_12 : std_logic;
  signal lbl1_cm_n_13, lbl1_cm_n_14, lbl1_cm_n_15, lbl1_cm_n_16, lbl1_cm_n_19 : std_logic;
  signal lbl1_cm_n_21, lbl1_cm_n_22, lbl1_cm_n_23, lbl1_cm_n_24, lbl1_cm_n_25 : std_logic;
  signal lbl1_cm_n_26, lbl1_cm_n_27, lbl1_cm_n_28, lbl1_cm_n_29, lbl1_cm_n_30 : std_logic;
  signal lbl1_cm_n_31, lbl1_cm_n_38, lbl1_cm_n_52, lbl1_cm_n_53, lbl1_cm_n_54 : std_logic;
  signal lbl1_cm_n_55, lbl1_cm_n_364_BAR, lbl1_cw_n_1, lbl1_cw_n_2, lbl1_cw_n_3 : std_logic;
  signal lbl1_cw_n_4, lbl1_cw_n_5, lbl1_cw_n_6, lbl1_cw_n_7, lbl1_cw_n_8 : std_logic;
  signal lbl1_cw_n_9, lbl1_cw_n_10, lbl1_cw_n_11, lbl1_cw_n_12, lbl1_cw_n_13 : std_logic;
  signal lbl1_cw_n_14, lbl1_cw_n_15, lbl1_cw_n_16, lbl1_cw_prev_incr, lbl1_cx_n_1 : std_logic;
  signal lbl1_cx_n_2, lbl1_cx_n_3, lbl1_cx_n_4, lbl1_cx_n_5, lbl1_cx_n_6 : std_logic;
  signal lbl1_cx_n_7, lbl1_cx_n_8, lbl1_cx_n_9, lbl1_cx_n_10, lbl1_cx_prev_incr : std_logic;
  signal lbl1_cy_n_1, lbl1_cy_n_2, lbl1_cy_n_3, lbl1_cy_n_4, lbl1_cy_n_5 : std_logic;
  signal lbl1_cy_n_6, lbl1_cy_n_7, lbl1_cy_n_8, lbl1_cy_n_9, lbl1_cy_n_10 : std_logic;
  signal lbl1_cy_prev_incr, lbl1_me_clr, lbl1_me_rw, lbl1_ready_clr, lbl1_ready_rw : std_logic;
  signal lbl1_rw_n_0, lbl1_rw_n_1, lbl1_rw_n_2, lbl1_rw_n_3, lbl1_rw_n_4 : std_logic;
  signal lbl1_rw_n_5, lbl1_rw_n_6, lbl1_rw_n_7, lbl1_rw_n_8, lbl1_rw_n_9 : std_logic;
  signal lbl1_rw_n_10, lbl1_rw_n_11, lbl1_rw_n_12, lbl1_rw_n_13, lbl1_rw_n_14 : std_logic;
  signal lbl1_rw_n_15, lbl1_rw_n_16, lbl1_rw_n_17, lbl1_rw_n_18, lbl1_rw_n_19 : std_logic;
  signal lbl1_rw_n_20, lbl1_rw_n_21, lbl1_rw_n_22, lbl1_rw_n_23, lbl1_rw_n_24 : std_logic;
  signal lbl1_rw_n_25, lbl1_rw_n_26, lbl1_rw_n_27, lbl1_rw_n_28, lbl1_rw_n_29 : std_logic;
  signal lbl1_rw_n_30, lbl1_rw_n_31, lbl1_rw_n_32, lbl1_rw_n_33, lbl1_rw_n_34 : std_logic;
  signal lbl1_rw_n_35, lbl1_rw_n_36, lbl1_rw_n_37, lbl1_rw_n_38, lbl1_rw_n_39 : std_logic;
  signal lbl1_rw_n_40, lbl1_rw_n_41, lbl1_rw_n_42, lbl1_rw_n_43, lbl1_rw_n_44 : std_logic;
  signal lbl1_rw_n_45, lbl1_rw_n_46, lbl1_rw_n_47, lbl1_rw_n_48, lbl1_rw_n_49 : std_logic;
  signal lbl1_rw_n_50, lbl1_rw_n_51, lbl1_rw_n_52, lbl1_rw_n_53, lbl1_rw_n_54 : std_logic;
  signal lbl1_rw_n_55, lbl1_rw_n_56, lbl1_rw_n_57, lbl1_rw_n_58, lbl1_rw_n_59 : std_logic;
  signal lbl1_rw_n_60, lbl1_rw_n_61, lbl1_rw_n_62, lbl1_rw_n_63, lbl1_rw_n_64 : std_logic;
  signal lbl1_rw_n_65, lbl1_rw_n_66, lbl1_rw_n_67, lbl1_rw_n_68, lbl1_rw_n_69 : std_logic;
  signal lbl1_rw_n_70, lbl1_rw_n_71, lbl1_rw_n_72, lbl1_rw_n_73, lbl1_rw_n_74 : std_logic;
  signal lbl1_rw_n_75, lbl1_rw_n_76, lbl1_rw_n_77, lbl1_rw_n_78, lbl1_rw_n_79 : std_logic;
  signal lbl1_rw_n_80, lbl1_rw_n_81, lbl1_rw_n_82, lbl1_rw_n_83, lbl1_rw_n_84 : std_logic;
  signal lbl1_rw_n_85, lbl1_rw_n_86, lbl1_rw_n_87, lbl1_rw_n_94, lbl1_rw_n_96 : std_logic;
  signal lbl1_rw_n_97, lbl1_rw_rst, lbl1_we_clr, lbl1_we_rw, lbl1_x_incr1 : std_logic;
  signal lbl1_x_incr2, lbl1_x_incr3, lbl1_y_incr1, lbl1_y_incr2, lbl1_y_incr3 : std_logic;
  signal lbl2_dec0_n_0, lbl2_dec0_n_1, lbl2_dec0_n_2, lbl2_dec0_n_3, lbl2_dec0_n_5 : std_logic;
  signal lbl2_dec1_n_0, lbl2_dec1_n_1, lbl2_dec1_n_2, lbl2_dec1_n_3, lbl2_dec1_n_5 : std_logic;
  signal lbl2_hscr_n_0, lbl2_hscr_n_1, lbl2_hscr_n_2, lbl2_hscr_n_6, lbl2_hscr_n_9 : std_logic;
  signal lbl2_hscr_n_10, lbl2_hscr_n_11, lbl2_hscr_n_12, lbl2_hscr_n_13, lbl2_hscr_n_14 : std_logic;
  signal lbl2_hscr_n_15, lbl2_hscr_n_16, lbl2_hscr_n_17, lbl2_hscr_n_18, lbl2_hscr_n_19 : std_logic;
  signal lbl2_hscr_n_20, lbl2_hscr_n_21, lbl2_hscr_n_22, lbl2_hscr_n_23, lbl2_hscr_n_24 : std_logic;
  signal lbl2_hscr_n_25, lbl2_hscr_n_26, lbl2_hscr_n_27, lbl2_hscr_n_28, lbl2_hscr_n_29 : std_logic;
  signal lbl2_hscr_n_30, lbl2_hscr_n_31, lbl2_hscr_n_32, lbl2_hscr_n_33, lbl2_hscr_n_34 : std_logic;
  signal lbl2_hscr_n_35, lbl2_hscr_n_36, lbl2_hscr_n_37, lbl2_hscr_n_38, lbl2_hscr_n_39 : std_logic;
  signal lbl2_hscr_n_40, lbl2_hscr_n_41, lbl2_hscr_n_42, lbl2_hscr_n_43, lbl2_hscr_n_44 : std_logic;
  signal lbl2_hscr_n_45, lbl2_hscr_n_46, lbl2_hscr_n_47, lbl2_hscr_n_48, lbl2_hscr_n_49 : std_logic;
  signal lbl2_hscr_n_50, lbl2_hscr_n_51, lbl2_hscr_n_52, lbl2_hscr_n_53, lbl2_hscr_n_54 : std_logic;
  signal lbl2_hscr_n_55, lbl2_hscr_n_56, lbl2_hscr_n_57, lbl2_hscr_n_58, lbl2_hscr_n_59 : std_logic;
  signal lbl2_hscr_n_60, lbl2_hscr_n_61, lbl2_hscr_n_62, lbl2_hscr_n_63, lbl2_hscr_n_64 : std_logic;
  signal lbl2_hscr_n_65, lbl2_hscr_n_66, lbl2_hscr_n_67, lbl2_hscr_n_68, lbl2_hscr_n_70 : std_logic;
  signal lbl2_hscr_n_71, lbl2_hscr_n_72, lbl2_hscr_n_73, lbl2_hscr_n_74, lbl2_hscr_n_76 : std_logic;
  signal lbl2_hscr_n_77, lbl2_hscr_n_78, lbl2_hscr_n_79, lbl2_hscr_n_80, lbl2_hscr_n_81 : std_logic;
  signal lbl2_hscr_n_82, lbl2_hscr_n_83, lbl2_hscr_n_84, lbl2_hscr_n_85, lbl2_hscr_n_86 : std_logic;
  signal lbl2_hscr_n_87, lbl2_hscr_n_88, lbl2_hscr_n_89, lbl2_hscr_n_90, lbl2_hscr_n_91 : std_logic;
  signal lbl2_hscr_n_92, lbl2_hscr_n_93, lbl2_hscr_n_94, lbl2_hscr_n_95, lbl2_hscr_n_96 : std_logic;
  signal lbl2_hscr_n_97, lbl2_hscr_n_98, lbl2_hscr_n_99, lbl2_hscr_n_100, lbl2_hscr_n_101 : std_logic;
  signal lbl2_hscr_n_102, lbl2_hscr_n_103, lbl2_hscr_n_104, lbl2_hscr_n_105, lbl2_hscr_n_106 : std_logic;
  signal lbl2_hscr_n_107, lbl2_hscr_n_108, lbl2_hscr_n_109, lbl2_hscr_n_110, lbl2_hscr_n_111 : std_logic;
  signal lbl2_hscr_n_112, lbl2_hscr_n_113, lbl2_hscr_n_114, lbl2_hscr_n_115, lbl2_hscr_n_116 : std_logic;
  signal lbl2_hscr_n_117, lbl2_hscr_n_118, lbl2_hscr_n_119, lbl2_hscr_n_120, lbl2_hscr_n_121 : std_logic;
  signal lbl2_hscr_n_122, lbl2_hscr_n_123, lbl2_hscr_n_124, lbl2_hscr_n_125, lbl2_hscr_n_126 : std_logic;
  signal lbl2_hscr_n_127, lbl2_hscr_n_128, lbl2_hscr_n_129, lbl2_hscr_n_130, lbl2_hscr_n_131 : std_logic;
  signal lbl2_hscr_n_132, lbl2_hscr_n_133, lbl2_hscr_n_134, lbl2_hscr_n_135, lbl2_hscr_n_136 : std_logic;
  signal lbl2_hscr_n_137, lbl2_hscr_n_138, lbl2_hscr_n_139, lbl2_hscr_n_140, lbl2_hscr_n_141 : std_logic;
  signal lbl2_hscr_n_142, lbl2_hscr_n_143, lbl2_hscr_n_144, lbl2_hscr_n_145, lbl2_hscr_n_146 : std_logic;
  signal lbl2_hscr_n_147, lbl2_hscr_n_148, lbl2_hscr_n_149, lbl2_hscr_n_150, lbl2_hscr_n_151 : std_logic;
  signal lbl2_hscr_n_153, lbl2_hscr_n_154, lbl2_hscr_n_155, lbl2_hscr_n_156, lbl2_hscr_n_157 : std_logic;
  signal lbl2_hscr_n_158, lbl2_hscr_n_159, lbl2_hscr_n_160, lbl2_hscr_n_161, lbl2_hscr_n_162 : std_logic;
  signal lbl2_hscr_n_163, lbl2_hscr_n_164, lbl2_hscr_n_165, lbl2_hscr_n_166, lbl2_hscr_n_167 : std_logic;
  signal lbl2_hscr_n_168, lbl2_hscr_n_169, lbl2_hscr_n_170, lbl2_hscr_n_171, lbl2_hscr_n_172 : std_logic;
  signal lbl2_hscr_n_173, lbl2_hscr_n_174, lbl2_hscr_n_175, lbl2_hscr_n_176, lbl2_hscr_n_177 : std_logic;
  signal lbl2_hscr_n_178, lbl2_hscr_n_179, lbl2_hscr_n_180, lbl2_hscr_n_181, lbl2_hscr_n_182 : std_logic;
  signal lbl2_hscr_n_183, lbl2_hscr_n_184, lbl2_hscr_n_185, lbl2_hscr_n_186, lbl2_hscr_n_187 : std_logic;
  signal lbl2_hscr_n_188, lbl2_hscr_n_189, lbl2_hscr_n_190, lbl2_hscr_n_191, lbl2_hscr_n_192 : std_logic;
  signal lbl2_hscr_n_193, lbl2_hscr_n_194, lbl2_hscr_n_195, lbl2_hscr_n_196, lbl2_hscr_n_197 : std_logic;
  signal lbl2_hscr_n_198, lbl2_hscr_n_199, lbl2_hscr_n_200, lbl2_hscr_n_201, lbl2_hscr_n_202 : std_logic;
  signal lbl2_hscr_n_203, lbl2_hscr_n_204, lbl2_hscr_n_205, lbl2_hscr_n_206, lbl2_hscr_n_207 : std_logic;
  signal lbl2_hscr_n_208, lbl2_hscr_n_209, lbl2_hscr_n_210, lbl2_hscr_n_211, lbl2_hscr_n_212 : std_logic;
  signal lbl2_hscr_n_213, lbl2_hscr_n_214, lbl2_hscr_n_215, lbl2_hscr_n_216, lbl2_hscr_n_217 : std_logic;
  signal lbl2_hscr_n_218, lbl2_hscr_n_219, lbl2_hscr_n_220, lbl2_hscr_n_221, lbl2_hscr_n_222 : std_logic;
  signal lbl2_hscr_n_223, lbl2_hscr_n_224, lbl2_hscr_n_225, lbl2_hscr_n_226, lbl2_hscr_n_227 : std_logic;
  signal lbl2_hscr_n_228, lbl2_hscr_n_229, lbl2_hscr_n_230, lbl2_hscr_n_231, lbl2_hscr_n_232 : std_logic;
  signal lbl2_hscr_n_233, lbl2_hscr_n_234, lbl2_hscr_n_235, lbl2_hscr_n_236, lbl2_hscr_n_237 : std_logic;
  signal lbl2_hscr_n_238, lbl2_hscr_n_239, lbl2_hscr_n_240, lbl2_hscr_n_241, lbl2_hscr_n_242 : std_logic;
  signal lbl2_hscr_n_243, lbl2_hscr_n_244, lbl2_hscr_n_245, lbl2_hscr_n_246, lbl2_hscr_n_247 : std_logic;
  signal lbl2_hscr_n_248, lbl2_hscr_n_249, lbl2_hscr_n_250, lbl2_hscr_n_251, lbl2_hscr_n_252 : std_logic;
  signal lbl2_hscr_n_253, lbl2_hscr_n_254, lbl2_hscr_n_255, lbl2_hscr_n_256, lbl2_hscr_n_257 : std_logic;
  signal lbl2_hscr_n_258, lbl2_hscr_n_259, lbl2_hscr_n_260, lbl2_hscr_n_261, lbl2_hscr_n_262 : std_logic;
  signal lbl2_hscr_n_263, lbl2_hscr_n_264, lbl2_hscr_n_265, lbl2_hscr_n_266, lbl2_hscr_n_267 : std_logic;
  signal lbl2_hscr_n_268, lbl2_hscr_n_269, lbl2_hscr_n_270, lbl2_hscr_n_271, lbl2_hscr_n_272 : std_logic;
  signal lbl2_hscr_n_273, lbl2_hscr_n_274, lbl2_hscr_n_275, lbl2_hscr_n_276, lbl2_hscr_n_277 : std_logic;
  signal lbl2_hscr_n_278, lbl2_hscr_n_279, lbl2_hscr_n_280, lbl2_hscr_n_281, lbl2_hscr_n_282 : std_logic;
  signal lbl2_hscr_n_283, lbl2_hscr_n_284, lbl2_hscr_n_285, lbl2_hscr_n_286, lbl2_hscr_n_287 : std_logic;
  signal lbl2_hscr_n_288, lbl2_hscr_n_289, lbl2_hscr_n_290, lbl2_hscr_n_291, lbl2_hscr_n_292 : std_logic;
  signal lbl2_hscr_n_293, lbl2_hscr_n_294, lbl2_hscr_n_295, lbl2_hscr_n_296, lbl2_hscr_n_297 : std_logic;
  signal lbl2_hscr_n_298, lbl2_hscr_n_299, lbl2_hscr_n_300, lbl2_hscr_n_301, lbl2_hscr_n_302 : std_logic;
  signal lbl2_hscr_n_303, lbl2_hscr_n_304, lbl2_hscr_n_305, lbl2_hscr_n_306, lbl2_hscr_n_307 : std_logic;
  signal lbl2_hscr_n_308, lbl2_hscr_n_309, lbl2_hscr_n_310, lbl2_hscr_n_311, lbl2_hscr_n_312 : std_logic;
  signal lbl2_hscr_n_313, lbl2_hscr_n_314, lbl2_hscr_n_315, lbl2_hscr_n_316, lbl2_hscr_n_317 : std_logic;
  signal lbl2_hscr_n_318, lbl2_hscr_n_319, lbl2_hscr_n_320, lbl2_hscr_n_321, lbl2_hscr_n_322 : std_logic;
  signal lbl2_hscr_n_323, lbl2_hscr_n_324, lbl2_hscr_n_325, lbl2_hscr_n_326, lbl2_hscr_n_327 : std_logic;
  signal lbl2_hscr_n_328, lbl2_hscr_n_329, lbl2_hscr_n_330, lbl2_hscr_n_331, lbl2_hscr_n_332 : std_logic;
  signal lbl2_hscr_n_333, lbl2_hscr_n_334, lbl2_hscr_n_335, lbl2_hscr_n_336, lbl2_hscr_n_337 : std_logic;
  signal lbl2_hscr_n_338, lbl2_hscr_n_339, lbl2_hscr_n_340, lbl2_hscr_n_341, lbl2_hscr_n_342 : std_logic;
  signal lbl2_hscr_n_343, lbl2_hscr_n_344, lbl2_hscr_n_345, lbl2_hscr_n_346, lbl2_hscr_n_347 : std_logic;
  signal lbl2_hscr_n_348, lbl2_hscr_n_349, lbl2_hscr_n_350, lbl2_hscr_n_351, lbl2_hscr_n_352 : std_logic;
  signal lbl2_hscr_n_353, lbl2_hscr_n_354, lbl2_hscr_n_355, lbl2_hscr_n_356, lbl2_hscr_n_357 : std_logic;
  signal lbl2_hscr_n_358, lbl2_hscr_n_359, lbl2_hscr_n_360, lbl2_hscr_n_361, lbl2_hscr_n_362 : std_logic;
  signal lbl2_hscr_n_363, lbl2_hscr_n_364, lbl2_hscr_n_365, lbl2_hscr_n_366, lbl2_hscr_n_367 : std_logic;
  signal lbl2_hscr_n_368, lbl2_hscr_n_369, lbl2_hscr_n_370, lbl2_hscr_n_371, lbl2_hscr_n_400 : std_logic;
  signal lbl2_hscr_n_401, lbl2_n_0, lbl2_n_1, lbl2_n_2, lbl2_n_3 : std_logic;
  signal lbl2_n_4, lbl2_n_5, lbl2_n_6, lbl2_n_7, lbl2_n_8 : std_logic;
  signal lbl2_n_9, lbl2_n_10, lbl2_n_11, lbl2_n_12, lbl2_n_13 : std_logic;
  signal lbl2_n_14, lbl2_n_15, lbl2_n_16, lbl2_n_17, lbl2_n_18 : std_logic;
  signal lbl2_n_19, lbl2_n_20, lbl2_n_21, lbl2_n_22, lbl2_n_23 : std_logic;
  signal lbl2_n_24, lbl2_n_25, lbl2_n_26, lbl2_n_27, lbl2_n_28 : std_logic;
  signal lbl2_n_29, lbl2_n_30, lbl2_n_31, lbl2_n_32, lbl2_n_33 : std_logic;
  signal lbl2_n_34, lbl2_n_35, lbl2_n_36, lbl2_n_37, lbl2_n_38 : std_logic;
  signal lbl2_n_39, lbl2_n_40, lbl2_n_41, lbl2_n_42, lbl2_n_43 : std_logic;
  signal lbl2_n_44, lbl2_n_45, lbl2_n_46, lbl2_n_47, lbl2_n_48 : std_logic;
  signal lbl2_n_49, lbl2_n_50, lbl2_n_51, lbl2_n_52, lbl2_n_53 : std_logic;
  signal lbl2_n_59, lbl2_n_60, lbl2_n_65, lbl2_n_66, lbl2_n_67 : std_logic;
  signal lbl2_n_68, lbl2_n_69, lbl2_n_70, lbl2_n_71, lbl2_n_72 : std_logic;
  signal lbl2_n_73, lbl2_n_74, lbl2_n_75, lbl2_n_77, lbl2_n_78 : std_logic;
  signal lbl2_n_79, lbl2_n_81, lbl2_n_82, lbl2_n_83, lbl2_n_84 : std_logic;
  signal lbl2_n_85, lbl2_n_86, lbl2_n_87, lbl2_n_88, lbl2_n_89 : std_logic;
  signal lbl2_n_90, lbl2_n_91, lbl2_n_92, lbl2_n_93, lbl2_n_94 : std_logic;
  signal lbl2_n_95, lbl2_n_96, lbl2_n_97, lbl2_n_98, lbl2_n_99 : std_logic;
  signal lbl2_n_100, lbl2_n_101, lbl2_n_102, lbl2_n_103, lbl2_n_104 : std_logic;
  signal lbl2_n_105, lbl2_n_106, lbl2_n_107, lbl2_n_108, lbl2_n_109 : std_logic;
  signal lbl2_n_110, lbl2_n_111, lbl2_n_113, lbl2_n_114, lbl2_n_115 : std_logic;
  signal lbl2_n_116, lbl2_n_117, lbl2_n_118, lbl2_n_119, lbl2_n_120 : std_logic;
  signal lbl2_n_122, lbl2_n_123, lbl2_n_124, lbl2_n_125, lbl2_n_126 : std_logic;
  signal lbl2_n_127, lbl2_n_128, lbl2_n_129, lbl2_n_130, lbl2_n_131 : std_logic;
  signal lbl2_n_132, lbl2_n_133, lbl2_n_134, lbl2_n_135, lbl2_n_136 : std_logic;
  signal lbl2_n_137, lbl2_n_138, lbl2_n_139, lbl2_n_140, lbl2_n_141 : std_logic;
  signal lbl2_n_142, lbl2_n_146, lbl2_n_147, lbl2_n_148, lbl2_n_149 : std_logic;
  signal lbl2_n_150, lbl2_n_151, lbl2_n_152, lbl2_n_153, lbl2_n_154 : std_logic;
  signal lbl2_n_156, lbl2_n_158, lbl2_n_189, lbl2_n_190, lbl2_n_227 : std_logic;
  signal lbl2_n_228, lbl2_n_229, lbl2_n_230, lbl2_pxl_n_0, lbl2_pxl_n_1 : std_logic;
  signal lbl2_pxl_n_2, lbl2_pxl_n_3, lbl2_pxl_n_5, lbl2_pxl_n_6, lbl2_pxl_n_7 : std_logic;
  signal lbl2_pxl_n_8, lbl2_pxl_n_9, lbl2_pxl_n_10, lbl2_pxl_n_11, lbl2_pxl_n_12 : std_logic;
  signal lbl2_pxl_n_13, lbl2_pxl_n_14, lbl2_pxl_n_15, lbl2_pxl_n_16, lbl2_pxl_n_17 : std_logic;
  signal lbl2_pxl_n_18, lbl2_pxl_n_19, lbl2_pxl_n_20, lbl2_pxl_n_21, lbl2_pxl_n_22 : std_logic;
  signal lbl2_pxl_n_23, lbl2_pxl_n_24, lbl2_pxl_n_25, lbl2_pxl_n_26, lbl2_pxl_n_27 : std_logic;
  signal lbl2_pxl_n_28, lbl2_pxl_n_29, lbl2_pxl_n_30, lbl2_pxl_n_31, lbl2_pxl_n_32 : std_logic;
  signal lbl2_pxl_n_33, lbl2_pxl_n_34, lbl2_pxl_n_35, lbl2_pxl_n_36, lbl2_pxl_n_37 : std_logic;
  signal lbl2_pxl_n_38, lbl2_pxl_n_39, lbl2_pxl_n_40, lbl2_pxl_n_41, lbl2_pxl_n_42 : std_logic;
  signal lbl2_pxl_n_43, lbl2_pxl_n_44, lbl2_pxl_n_45, lbl2_pxl_n_46, lbl2_pxl_n_47 : std_logic;
  signal lbl2_pxl_n_48, lbl2_pxl_n_49, lbl2_pxl_n_50, lbl2_pxl_n_51, lbl2_pxl_n_52 : std_logic;
  signal lbl2_pxl_n_53, lbl2_pxl_n_54, lbl2_pxl_n_55, lbl2_pxl_n_56, lbl2_pxl_n_57 : std_logic;
  signal lbl2_pxl_n_58, lbl2_pxl_n_59, lbl2_pxl_n_60, lbl2_pxl_n_61, lbl2_pxl_n_62 : std_logic;
  signal lbl2_pxl_n_63, lbl2_pxl_n_64, lbl2_pxl_n_65, lbl2_pxl_n_66, lbl2_pxl_n_67 : std_logic;
  signal lbl2_pxl_n_68, lbl2_pxl_n_69, lbl2_pxl_n_70, lbl2_pxl_n_71, lbl2_pxl_n_72 : std_logic;
  signal lbl2_pxl_n_73, lbl2_pxl_n_74, lbl2_pxl_n_75, lbl2_pxl_n_76, lbl2_pxl_n_77 : std_logic;
  signal lbl2_pxl_n_78, lbl2_pxl_n_79, lbl2_pxl_n_80, lbl2_pxl_n_81, lbl2_pxl_n_82 : std_logic;
  signal lbl2_pxl_n_83, lbl2_pxl_n_84, lbl2_pxl_n_85, lbl2_pxl_n_86, lbl2_pxl_n_87 : std_logic;
  signal lbl2_pxl_n_88, lbl2_pxl_n_89, lbl2_pxl_n_90, lbl2_pxl_n_91, lbl2_pxl_n_92 : std_logic;
  signal lbl2_pxl_n_93, lbl2_pxl_n_94, lbl2_pxl_n_95, lbl2_pxl_n_96, lbl2_pxl_n_97 : std_logic;
  signal lbl2_pxl_n_98, lbl2_pxl_n_99, lbl2_pxl_n_100, lbl2_pxl_n_101, lbl2_pxl_n_102 : std_logic;
  signal lbl2_pxl_n_103, lbl2_pxl_n_104, lbl2_pxl_n_105, lbl2_pxl_n_106, lbl2_pxl_n_107 : std_logic;
  signal lbl2_pxl_n_108, lbl2_pxl_n_109, lbl2_pxl_n_110, lbl2_pxl_n_111, lbl2_pxl_n_112 : std_logic;
  signal lbl2_pxl_n_113, lbl2_pxl_n_114, lbl2_pxl_n_115, lbl2_pxl_n_116, lbl2_pxl_n_117 : std_logic;
  signal lbl2_pxl_n_118, lbl2_pxl_n_119, lbl2_pxl_n_120, lbl2_pxl_n_121, lbl2_pxl_n_122 : std_logic;
  signal lbl2_pxl_n_123, lbl2_pxl_n_124, lbl2_pxl_n_125, lbl2_pxl_n_126, lbl2_pxl_n_127 : std_logic;
  signal lbl2_pxl_n_128, lbl2_pxl_n_129, lbl2_pxl_n_130, lbl2_pxl_n_131, lbl2_pxl_n_132 : std_logic;
  signal lbl2_pxl_n_133, lbl2_pxl_n_134, lbl2_pxl_n_135, lbl2_pxl_n_136, lbl2_pxl_n_137 : std_logic;
  signal lbl2_pxl_n_138, lbl2_pxl_n_139, lbl2_pxl_n_140, lbl2_pxl_n_141, lbl2_pxl_n_142 : std_logic;
  signal lbl2_pxl_n_143, lbl2_pxl_n_144, lbl2_pxl_n_145, lbl2_pxl_n_146, lbl2_pxl_n_147 : std_logic;
  signal lbl2_pxl_n_148, lbl2_pxl_n_149, lbl2_pxl_n_150, lbl2_pxl_n_151, lbl2_pxl_n_152 : std_logic;
  signal lbl2_pxl_n_153, lbl2_pxl_n_154, lbl2_pxl_n_155, lbl2_pxl_n_156, lbl2_pxl_n_157 : std_logic;
  signal lbl2_pxl_n_158, lbl2_pxl_n_159, lbl2_pxl_n_160, lbl2_pxl_n_161, lbl2_pxl_n_162 : std_logic;
  signal lbl2_pxl_n_163, lbl2_pxl_n_164, lbl2_pxl_n_165, lbl2_pxl_n_166, lbl2_pxl_n_167 : std_logic;
  signal lbl2_pxl_n_168, lbl2_pxl_n_169, lbl2_pxl_n_170, lbl2_pxl_n_171, lbl2_pxl_n_172 : std_logic;
  signal lbl2_pxl_n_173, lbl2_pxl_n_174, lbl2_pxl_n_175, lbl2_pxl_n_176, lbl2_pxl_n_177 : std_logic;
  signal lbl2_pxl_n_178, lbl2_pxl_n_179, lbl2_pxl_n_180, lbl2_pxl_n_181, lbl2_pxl_n_182 : std_logic;
  signal lbl2_pxl_n_183, lbl2_pxl_n_184, lbl2_pxl_n_185, lbl2_pxl_n_186, lbl2_pxl_n_187 : std_logic;
  signal lbl2_pxl_n_188, lbl2_pxl_n_189, lbl2_pxl_n_190, lbl2_pxl_n_191, lbl2_pxl_n_192 : std_logic;
  signal lbl2_pxl_n_193, lbl2_pxl_n_194, lbl2_pxl_n_195, lbl2_pxl_n_196, lbl2_pxl_n_197 : std_logic;
  signal lbl2_pxl_n_198, lbl2_pxl_n_199, lbl2_pxl_n_200, lbl2_pxl_n_201, lbl2_pxl_n_202 : std_logic;
  signal lbl2_pxl_n_203, lbl2_pxl_n_205, lbl2_pxl_n_206, lbl2_pxl_n_207, lbl2_pxl_n_208 : std_logic;
  signal lbl2_pxl_n_210, lbl2_sdb_n_0, lbl2_sdb_n_1, lbl2_sdb_n_2, lbl2_sdb_n_3 : std_logic;
  signal lbl2_sdb_n_8, lbl2_sdb_n_9, lbl2_sdb_n_10, lbl2_sdb_n_11, lbl2_sdb_n_12 : std_logic;
  signal lbl2_sdb_n_13, lbl2_sdb_n_14, lbl2_sdb_n_15, lbl2_sdb_n_16, lbl2_sdb_n_17 : std_logic;
  signal lbl2_sdb_n_18, lbl2_sdb_n_19, lbl2_sdb_n_20, lbl2_sdb_n_21, lbl2_sdb_n_22 : std_logic;
  signal lbl2_sdb_n_23, lbl2_sdb_n_24, lbl2_sdb_n_25, lbl2_sdb_n_26, lbl2_sdb_n_27 : std_logic;
  signal lbl2_sdb_n_28, lbl2_sdb_n_29, lbl2_sdb_n_30, lbl2_sdb_n_31, lbl2_sdb_n_32 : std_logic;
  signal lbl2_sdb_n_33, lbl2_sdb_n_34, lbl2_sdb_n_35, lbl2_sdb_n_36, lbl2_sdb_n_37 : std_logic;
  signal lbl2_sdb_n_38, lbl2_sdb_n_39, lbl2_sdb_n_40, lbl2_sdb_n_41, lbl2_sdb_n_42 : std_logic;
  signal lbl2_sdb_n_43, lbl2_sdb_n_44, lbl2_sdb_n_45, lbl2_sdb_n_46, lbl2_sdb_n_47 : std_logic;
  signal lbl2_sdb_n_48, lbl2_sdb_n_49, lbl2_sdb_n_50, lbl2_sdb_n_51, lbl2_sdb_n_52 : std_logic;
  signal lbl2_sdb_n_53, lbl2_sdb_n_54, lbl2_sdb_n_55, lbl2_sdb_n_56, lbl2_sdb_n_57 : std_logic;
  signal lbl2_sdb_n_58, lbl2_sdb_n_59, lbl2_sdb_n_60, lbl2_sdb_n_61, lbl2_sdb_n_62 : std_logic;
  signal lbl2_sdb_n_63, lbl2_sdb_n_64, lbl2_sdb_n_65, lbl2_sdb_n_66, lbl2_sdb_n_67 : std_logic;
  signal lbl2_sdb_n_68, lbl2_sdb_n_70, lbl2_sdb_n_71, lbl2_sdb_n_72, lbl2_sdb_n_73 : std_logic;
  signal lbl2_sdb_n_74, lbl2_sdb_n_75, lbl2_sdb_n_76, lbl2_sdb_n_77, lbl2_sdb_n_78 : std_logic;
  signal lbl2_sdb_n_79, lbl2_sdb_n_80, lbl2_sdb_n_81, lbl2_sdb_n_82, lbl2_sdb_n_83 : std_logic;
  signal lbl2_sdb_n_85, lbl2_sdb_n_86, lbl2_sdb_n_87, lbl2_sdb_n_88, lbl2_sdb_n_89 : std_logic;
  signal lbl2_sdb_n_90, lbl2_sdb_n_91, lbl2_sdb_n_92, lbl2_sdb_n_93, lbl2_sdb_n_94 : std_logic;
  signal lbl2_sdb_n_95, lbl2_sdb_n_96, lbl2_sdb_n_97, lbl2_sdb_n_98, lbl2_sdb_n_99 : std_logic;
  signal lbl2_sdb_n_100, lbl2_sdb_n_101, lbl2_sdb_n_102, lbl2_sdb_n_103, lbl2_sdb_n_104 : std_logic;
  signal lbl2_sdb_n_105, lbl2_sdb_n_106, lbl2_sdb_n_107, lbl2_sdb_n_108, lbl2_sdb_n_109 : std_logic;
  signal lbl2_sdb_n_110, lbl2_sdb_n_111, lbl2_sdb_n_112, lbl2_sdb_n_113, lbl2_sdb_n_114 : std_logic;
  signal lbl2_sdb_n_115, lbl2_sdb_n_116, lbl2_sdb_n_117, lbl2_sdb_n_118, lbl2_sdb_n_119 : std_logic;
  signal lbl2_sdb_n_120, lbl2_sdb_n_121, lbl2_sdb_n_122, lbl2_sdb_n_123, lbl2_sdb_n_124 : std_logic;
  signal lbl2_sdb_n_125, lbl2_sdb_n_126, lbl2_sdb_n_127, lbl2_sdb_n_128, lbl2_sdb_n_129 : std_logic;
  signal lbl2_sdb_n_130, lbl2_sdb_n_131, lbl2_sdb_n_132, lbl2_sdb_n_133, lbl2_sdb_n_134 : std_logic;
  signal lbl2_sdb_n_135, lbl2_sdb_n_136, lbl2_sdb_n_137, lbl2_sdb_n_138, lbl2_sdb_n_139 : std_logic;
  signal lbl2_sdb_n_140, lbl2_sdb_n_141, lbl2_sdb_n_142, lbl2_sdb_n_143, lbl2_sdb_n_144 : std_logic;
  signal lbl2_sdb_n_145, lbl2_sdb_n_146, lbl2_sdb_n_147, lbl2_sdb_n_148, lbl2_sdb_n_149 : std_logic;
  signal lbl2_sdb_n_150, lbl2_sdb_n_151, lbl2_sdb_n_152, lbl2_sdb_n_153, lbl2_sdb_n_154 : std_logic;
  signal lbl2_sdb_n_155, lbl2_sdb_n_156, lbl2_sdb_n_157, lbl2_sdb_n_158, lbl2_sdb_n_159 : std_logic;
  signal lbl2_sdb_n_160, lbl2_sdb_n_161, lbl2_sdb_n_162, lbl2_sdb_n_163, lbl2_sdb_n_164 : std_logic;
  signal lbl2_sdb_n_165, lbl2_sdb_n_166, lbl2_sdb_n_167, lbl2_sdb_n_168, lbl2_sdb_n_169 : std_logic;
  signal lbl2_sdb_n_170, lbl2_sdb_n_171, lbl2_sdb_n_172, lbl2_sdb_n_173, lbl2_sdb_n_174 : std_logic;
  signal lbl2_sdb_n_175, lbl2_sdb_n_176, lbl2_sdb_n_177, lbl2_sdb_n_178, lbl2_sdb_n_179 : std_logic;
  signal lbl2_sdb_n_180, lbl2_sdb_n_181, lbl2_sdb_n_182, lbl2_sdb_n_183, lbl2_sdb_n_184 : std_logic;
  signal lbl2_sdb_n_185, lbl2_sdb_n_186, lbl2_sdb_n_187, lbl2_sdb_n_188, lbl2_sdb_n_189 : std_logic;
  signal lbl2_sdb_n_190, lbl2_sdb_n_191, lbl2_sdb_n_192, lbl2_sdb_n_193, lbl2_sdb_n_194 : std_logic;
  signal lbl2_sdb_n_214, lbl3_temp2, lbl4_n_2, lbl4_n_3, lbl4_n_4 : std_logic;
  signal lbl4_n_5, lbl4_n_6, lbl4_n_7, lbl4_n_8, lbl4_n_9 : std_logic;
  signal lbl4_n_10, lbl4_n_12, lbl4_n_13, lbl4_n_14, lbl4_n_15 : std_logic;
  signal lbl4_n_16, lbl4_n_17, lbl4_n_18, lbl4_n_19, lbl4_n_20 : std_logic;
  signal lbl4_n_21, lbl4_n_22, lbl4_n_23, lbl4_n_24, lbl4_n_27 : std_logic;
  signal lbl4_n_28, lbl4_n_29, lbl4_n_30, lbl4_n_31, lbl4_n_32 : std_logic;
  signal lbl4_n_33, lbl4_n_34, lbl4_n_35, lbl4_n_36, lbl4_n_37 : std_logic;
  signal lbl4_n_38, lbl4_n_39, lbl4_n_41, lbl4_n_42, lbl4_n_43 : std_logic;
  signal lbl4_n_44, lbl4_n_45, lbl4_n_46, lbl4_n_47, lbl4_n_48 : std_logic;
  signal lbl4_n_49, lbl4_n_50, lbl4_n_51, lbl4_n_52, lbl4_n_53 : std_logic;
  signal lbl4_n_54, lbl4_n_55, lbl4_n_56, lbl4_n_57, lbl4_n_58 : std_logic;
  signal lbl4_n_59, lbl4_n_60, lbl4_n_61, lbl4_n_62, lbl4_n_63 : std_logic;
  signal lbl4_n_64, lbl4_n_65, lbl4_n_66, lbl4_n_67, lbl4_n_68 : std_logic;
  signal lbl4_n_69, lbl4_n_70, lbl4_n_71, lbl4_n_72, lbl4_n_73 : std_logic;
  signal lbl4_n_74, lbl4_n_75, lbl4_n_76, lbl4_n_77, lbl4_n_78 : std_logic;
  signal lbl4_n_79, lbl4_n_80, lbl4_n_81, lbl4_n_82, lbl4_n_83 : std_logic;
  signal lbl4_n_84, lbl4_n_85, lbl4_n_86, lbl4_n_87, lbl4_n_88 : std_logic;
  signal lbl4_n_89, lbl4_n_90, lbl4_n_91, lbl4_n_92, lbl4_n_93 : std_logic;
  signal lbl4_n_94, lbl4_n_95, lbl4_n_96, lbl4_n_97, lbl4_n_98 : std_logic;
  signal lbl4_n_99, lbl4_n_100, lbl4_n_101, lbl4_n_102, lbl4_n_103 : std_logic;
  signal lbl4_n_104, lbl4_n_105, lbl4_n_106, lbl4_n_107, lbl4_n_108 : std_logic;
  signal lbl4_n_109, lbl4_n_110, lbl4_n_111, lbl4_n_112, lbl4_n_113 : std_logic;
  signal lbl4_n_114, lbl4_n_115, lbl4_n_116, lbl4_n_117, lbl4_n_118 : std_logic;
  signal lbl4_n_119, lbl4_n_120, lbl4_n_121, lbl4_n_122, lbl4_n_123 : std_logic;
  signal lbl4_n_124, lbl4_n_125, lbl4_n_126, lbl4_n_127, lbl4_n_130 : std_logic;
  signal lbl4_n_134, lbl4_n_137, lbl4_n_138, lbl4_n_140, lbl4_n_141 : std_logic;
  signal lbl4_n_142, lbl4_n_147, lbl5_beep_en, lbl5_crash_en, lbl5_en0_csa_tree_lt_140_15_groupi_n_0 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_2, lbl5_en0_csa_tree_lt_140_15_groupi_n_3, lbl5_en0_csa_tree_lt_140_15_groupi_n_4, lbl5_en0_csa_tree_lt_140_15_groupi_n_5, lbl5_en0_csa_tree_lt_140_15_groupi_n_6 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_7, lbl5_en0_csa_tree_lt_140_15_groupi_n_8, lbl5_en0_csa_tree_lt_140_15_groupi_n_9, lbl5_en0_csa_tree_lt_140_15_groupi_n_10, lbl5_en0_csa_tree_lt_140_15_groupi_n_11 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_12, lbl5_en0_csa_tree_lt_140_15_groupi_n_13, lbl5_en0_csa_tree_lt_140_15_groupi_n_14, lbl5_en0_csa_tree_lt_140_15_groupi_n_15, lbl5_en0_csa_tree_lt_140_15_groupi_n_16 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_17, lbl5_en0_csa_tree_lt_140_15_groupi_n_18, lbl5_en0_csa_tree_lt_140_15_groupi_n_19, lbl5_en0_csa_tree_lt_140_15_groupi_n_20, lbl5_en0_csa_tree_lt_140_15_groupi_n_21 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_22, lbl5_en0_csa_tree_lt_140_15_groupi_n_23, lbl5_en0_csa_tree_lt_140_15_groupi_n_24, lbl5_en0_csa_tree_lt_140_15_groupi_n_25, lbl5_en0_csa_tree_lt_140_15_groupi_n_26 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_27, lbl5_en0_csa_tree_lt_140_15_groupi_n_28, lbl5_en0_csa_tree_lt_140_15_groupi_n_29, lbl5_en0_csa_tree_lt_140_15_groupi_n_30, lbl5_en0_csa_tree_lt_140_15_groupi_n_31 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_32, lbl5_en0_csa_tree_lt_140_15_groupi_n_33, lbl5_en0_csa_tree_lt_140_15_groupi_n_34, lbl5_en0_csa_tree_lt_140_15_groupi_n_36, lbl5_en0_csa_tree_lt_140_15_groupi_n_37 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_38, lbl5_en0_csa_tree_lt_140_15_groupi_n_39, lbl5_en0_csa_tree_lt_140_15_groupi_n_40, lbl5_en0_csa_tree_lt_140_15_groupi_n_41, lbl5_en0_csa_tree_lt_140_15_groupi_n_42 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_43, lbl5_en0_csa_tree_lt_140_15_groupi_n_44, lbl5_en0_csa_tree_lt_140_15_groupi_n_45, lbl5_en0_csa_tree_lt_140_15_groupi_n_46, lbl5_en0_csa_tree_lt_140_15_groupi_n_47 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_48, lbl5_en0_csa_tree_lt_140_15_groupi_n_49, lbl5_en0_csa_tree_lt_140_15_groupi_n_50, lbl5_en0_csa_tree_lt_140_15_groupi_n_51, lbl5_en0_csa_tree_lt_140_15_groupi_n_52 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_53, lbl5_en0_csa_tree_lt_140_15_groupi_n_54, lbl5_en0_csa_tree_lt_140_15_groupi_n_55, lbl5_en0_csa_tree_lt_140_15_groupi_n_56, lbl5_en0_csa_tree_lt_140_15_groupi_n_57 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_58, lbl5_en0_csa_tree_lt_140_15_groupi_n_59, lbl5_en0_csa_tree_lt_140_15_groupi_n_60, lbl5_en0_csa_tree_lt_140_15_groupi_n_61, lbl5_en0_csa_tree_lt_140_15_groupi_n_62 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_63, lbl5_en0_csa_tree_lt_140_15_groupi_n_64, lbl5_en0_csa_tree_lt_140_15_groupi_n_65, lbl5_en0_csa_tree_lt_140_15_groupi_n_66, lbl5_en0_csa_tree_lt_140_15_groupi_n_67 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_68, lbl5_en0_csa_tree_lt_140_15_groupi_n_69, lbl5_en0_csa_tree_lt_140_15_groupi_n_112, lbl5_en0_csa_tree_lt_140_15_groupi_n_114, lbl5_en0_csa_tree_lt_140_15_groupi_n_118 : std_logic;
  signal lbl5_en0_csa_tree_lt_140_15_groupi_n_119, lbl5_en0_csa_tree_lt_140_15_groupi_n_120, lbl5_en0_csa_tree_lt_140_15_groupi_n_121, lbl5_en0_csa_tree_lt_140_15_groupi_n_123, lbl5_en0_csa_tree_lt_140_15_groupi_n_124 : std_logic;
  signal lbl5_en0_frozen_boost, lbl5_en0_inc_add_127_23_n_0, lbl5_en0_inc_add_127_23_n_2, lbl5_en0_inc_add_127_23_n_4, lbl5_en0_inc_add_127_23_n_6 : std_logic;
  signal lbl5_en0_inc_add_127_23_n_8, lbl5_en0_inc_add_127_23_n_10, lbl5_en0_inc_add_127_23_n_12, lbl5_en0_inc_add_127_23_n_14, lbl5_en0_inc_add_127_23_n_16 : std_logic;
  signal lbl5_en0_inc_add_127_23_n_18, lbl5_en0_inc_add_127_23_n_20, lbl5_en0_inc_add_127_23_n_22, lbl5_en0_inc_add_127_23_n_24, lbl5_en0_inc_add_127_23_n_26 : std_logic;
  signal lbl5_en0_inc_add_127_23_n_28, lbl5_en0_inc_add_127_23_n_30, lbl5_en0_inc_add_127_23_n_32, lbl5_en0_n_0, lbl5_en0_n_1 : std_logic;
  signal lbl5_en0_n_2, lbl5_en0_n_3, lbl5_en0_n_4, lbl5_en0_n_5, lbl5_en0_n_6 : std_logic;
  signal lbl5_en0_n_7, lbl5_en0_n_8, lbl5_en0_n_9, lbl5_en0_n_10, lbl5_en0_n_11 : std_logic;
  signal lbl5_en0_n_12, lbl5_en0_n_13, lbl5_en0_n_14, lbl5_en0_n_15, lbl5_en0_n_16 : std_logic;
  signal lbl5_en0_n_17, lbl5_en0_n_18, lbl5_en0_n_19, lbl5_en0_n_20, lbl5_en0_n_21 : std_logic;
  signal lbl5_en0_n_22, lbl5_en0_n_23, lbl5_en0_n_24, lbl5_en0_n_25, lbl5_en0_n_26 : std_logic;
  signal lbl5_en0_n_27, lbl5_en0_n_28, lbl5_en0_n_29, lbl5_en0_n_30, lbl5_en0_n_31 : std_logic;
  signal lbl5_en0_n_32, lbl5_en0_n_33, lbl5_en0_n_34, lbl5_en0_n_35, lbl5_en0_n_36 : std_logic;
  signal lbl5_en0_n_37, lbl5_en0_n_38, lbl5_en0_n_39, lbl5_en0_n_40, lbl5_en0_n_41 : std_logic;
  signal lbl5_en0_n_42, lbl5_en0_n_43, lbl5_en0_n_44, lbl5_en0_n_45, lbl5_en0_n_46 : std_logic;
  signal lbl5_en0_n_47, lbl5_en0_n_48, lbl5_en0_n_49, lbl5_en0_n_50, lbl5_en0_n_51 : std_logic;
  signal lbl5_en0_n_52, lbl5_en0_n_53, lbl5_en0_n_54, lbl5_en0_n_55, lbl5_en0_n_56 : std_logic;
  signal lbl5_en0_n_57, lbl5_en0_n_58, lbl5_en0_n_59, lbl5_en0_n_60, lbl5_en0_n_61 : std_logic;
  signal lbl5_en0_n_62, lbl5_en0_n_63, lbl5_en0_n_64, lbl5_en0_n_65, lbl5_en0_n_66 : std_logic;
  signal lbl5_en0_n_67, lbl5_en0_n_68, lbl5_en0_n_69, lbl5_en0_n_70, lbl5_en0_n_71 : std_logic;
  signal lbl5_en0_n_72, lbl5_en0_n_73, lbl5_en0_n_74, lbl5_en0_n_75, lbl5_en0_n_76 : std_logic;
  signal lbl5_en0_n_77, lbl5_en0_n_78, lbl5_en0_n_79, lbl5_en0_n_80, lbl5_en0_n_81 : std_logic;
  signal lbl5_en0_n_82, lbl5_en0_n_83, lbl5_en0_n_84, lbl5_en0_n_85, lbl5_en0_n_86 : std_logic;
  signal lbl5_en0_n_87, lbl5_en0_n_88, lbl5_en0_n_89, lbl5_en0_n_90, lbl5_en0_n_91 : std_logic;
  signal lbl5_en0_n_92, lbl5_en0_n_93, lbl5_en0_n_94, lbl5_en0_n_95, lbl5_en0_n_96 : std_logic;
  signal lbl5_en0_n_97, lbl5_en0_n_98, lbl5_en0_n_99, lbl5_en0_n_100, lbl5_en0_n_101 : std_logic;
  signal lbl5_en0_n_102, lbl5_en0_n_103, lbl5_en0_n_104, lbl5_en0_n_105, lbl5_en0_n_106 : std_logic;
  signal lbl5_en0_n_107, lbl5_en0_n_108, lbl5_en0_n_109, lbl5_en0_n_110, lbl5_en0_n_111 : std_logic;
  signal lbl5_en0_n_112, lbl5_en0_n_113, lbl5_en0_n_114, lbl5_en0_n_115, lbl5_en0_n_116 : std_logic;
  signal lbl5_en0_n_117, lbl5_en0_n_118, lbl5_en0_n_119, lbl5_en0_n_120, lbl5_en0_n_121 : std_logic;
  signal lbl5_en0_n_122, lbl5_en0_n_123, lbl5_en0_n_124, lbl5_en0_n_125, lbl5_en0_n_126 : std_logic;
  signal lbl5_en0_n_127, lbl5_en0_n_128, lbl5_en0_n_129, lbl5_en0_n_130, lbl5_en0_n_131 : std_logic;
  signal lbl5_en0_n_132, lbl5_en0_n_133, lbl5_en0_n_134, lbl5_en0_n_135, lbl5_en0_n_136 : std_logic;
  signal lbl5_en0_n_137, lbl5_en0_n_138, lbl5_en0_n_139, lbl5_en0_n_140, lbl5_en0_n_141 : std_logic;
  signal lbl5_en0_n_142, lbl5_en0_n_143, lbl5_en0_n_144, lbl5_en0_n_145, lbl5_en0_n_146 : std_logic;
  signal lbl5_en0_n_147, lbl5_en0_n_148, lbl5_en0_n_149, lbl5_en0_n_150, lbl5_en0_n_151 : std_logic;
  signal lbl5_en0_n_152, lbl5_en0_n_153, lbl5_en0_n_154, lbl5_en0_n_155, lbl5_en0_n_156 : std_logic;
  signal lbl5_en0_n_157, lbl5_en0_n_158, lbl5_en0_n_159, lbl5_en0_n_160, lbl5_en0_n_161 : std_logic;
  signal lbl5_en0_n_162, lbl5_en0_n_163, lbl5_en0_n_164, lbl5_en0_n_165, lbl5_en0_n_166 : std_logic;
  signal lbl5_en0_n_167, lbl5_en0_n_168, lbl5_en0_n_169, lbl5_en0_n_170, lbl5_en0_n_171 : std_logic;
  signal lbl5_en0_n_172, lbl5_en0_n_173, lbl5_en0_n_174, lbl5_en0_n_175, lbl5_en0_n_176 : std_logic;
  signal lbl5_en0_n_177, lbl5_en0_n_178, lbl5_en0_n_179, lbl5_en0_n_182, lbl5_en0_n_186 : std_logic;
  signal lbl5_en0_n_187, lbl5_en0_n_188, lbl5_en0_n_190, lbl5_en0_n_191, lbl5_en0_n_193 : std_logic;
  signal lbl5_en0_n_196, lbl5_en0_n_198, lbl5_en0_n_199, lbl5_en0_n_200, lbl5_en0_n_201 : std_logic;
  signal lbl5_en0_n_202, lbl5_en0_n_203, lbl5_en0_n_204, lbl5_en0_n_205, lbl5_en0_n_206 : std_logic;
  signal lbl5_en0_n_207, lbl5_en0_n_208, lbl5_en0_n_209, lbl5_en0_n_210, lbl5_en0_n_211 : std_logic;
  signal lbl5_en0_n_212, lbl5_en0_n_213, lbl5_en0_n_214, lbl5_en0_n_215, lbl5_en0_n_216 : std_logic;
  signal lbl5_en0_n_218, lbl5_en0_n_219, lbl5_en0_n_220, lbl5_en0_n_221, lbl5_en0_n_222 : std_logic;
  signal lbl5_en0_n_223, lbl5_en0_n_224, lbl5_en0_n_225, lbl5_en0_n_226, lbl5_en0_n_227 : std_logic;
  signal lbl5_en0_n_228, lbl5_en0_n_229, lbl5_en0_n_230, lbl5_en0_n_231, lbl5_en0_n_232 : std_logic;
  signal lbl5_en0_n_233, lbl5_en0_n_234, lbl5_en0_n_235, lbl5_en0_n_236, lbl5_en0_n_237 : std_logic;
  signal lbl5_en0_n_238, lbl5_en0_n_239, lbl5_en0_n_240, lbl5_en0_n_241, lbl5_en0_n_242 : std_logic;
  signal lbl5_en0_n_243, lbl5_en0_n_244, lbl5_en0_n_245, lbl5_en0_n_246, lbl5_en0_n_247 : std_logic;
  signal lbl5_en0_n_248, lbl5_en0_n_249, lbl5_en0_n_250, lbl5_en0_n_251, lbl5_en0_n_252 : std_logic;
  signal lbl5_en0_n_253, lbl5_en0_n_254, lbl5_en0_n_255, lbl5_en0_n_256, lbl5_en0_n_257 : std_logic;
  signal lbl5_en0_n_258, lbl5_en0_n_259, lbl5_en0_n_260, lbl5_en0_n_261, lbl5_en0_n_263 : std_logic;
  signal lbl5_en0_n_264, lbl5_en0_n_265, lbl5_en0_n_266, lbl5_en0_n_267, lbl5_en0_n_268 : std_logic;
  signal lbl5_en0_n_269, lbl5_en0_n_270, lbl5_en0_n_271, lbl5_en0_n_272, lbl5_en0_n_273 : std_logic;
  signal lbl5_en0_n_274, lbl5_en0_n_276, lbl5_en0_n_277, lbl5_en0_n_278, lbl5_en0_n_280 : std_logic;
  signal lbl5_en0_n_281, lbl5_en0_n_282, lbl5_en0_n_283, lbl5_en0_n_284, lbl5_en0_n_285 : std_logic;
  signal lbl5_en0_n_286, lbl5_en0_n_287, lbl5_en0_n_288, lbl5_en0_n_289, lbl5_en0_n_290 : std_logic;
  signal lbl5_en0_n_291, lbl5_en0_n_292, lbl5_en0_n_293, lbl5_en0_n_294, lbl5_en0_n_295 : std_logic;
  signal lbl5_en0_n_296, lbl5_en0_n_297, lbl5_en0_n_298, lbl5_en0_n_299, lbl5_en0_n_300 : std_logic;
  signal lbl5_en0_n_301, lbl5_en0_n_302, lbl5_en0_n_303, lbl5_en0_n_304, lbl5_en0_n_305 : std_logic;
  signal lbl5_en0_n_306, lbl5_en0_n_307, lbl5_en0_n_308, lbl5_en0_n_309, lbl5_en0_n_310 : std_logic;
  signal lbl5_en0_n_311, lbl5_en0_n_312, lbl5_en0_n_313, lbl5_en0_n_314, lbl5_en0_n_315 : std_logic;
  signal lbl5_en0_n_316, lbl5_en0_n_327, lbl5_en0_n_328, lbl5_en0_n_329, lbl5_en0_prev_crash : std_logic;
  signal lbl5_en0_prev_engine, lbl5_en0_rst, lbl5_en1_csa_tree_lt_140_15_groupi_n_0, lbl5_en1_csa_tree_lt_140_15_groupi_n_2, lbl5_en1_csa_tree_lt_140_15_groupi_n_3 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_4, lbl5_en1_csa_tree_lt_140_15_groupi_n_5, lbl5_en1_csa_tree_lt_140_15_groupi_n_6, lbl5_en1_csa_tree_lt_140_15_groupi_n_7, lbl5_en1_csa_tree_lt_140_15_groupi_n_8 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_9, lbl5_en1_csa_tree_lt_140_15_groupi_n_10, lbl5_en1_csa_tree_lt_140_15_groupi_n_11, lbl5_en1_csa_tree_lt_140_15_groupi_n_12, lbl5_en1_csa_tree_lt_140_15_groupi_n_13 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_14, lbl5_en1_csa_tree_lt_140_15_groupi_n_15, lbl5_en1_csa_tree_lt_140_15_groupi_n_16, lbl5_en1_csa_tree_lt_140_15_groupi_n_17, lbl5_en1_csa_tree_lt_140_15_groupi_n_18 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_19, lbl5_en1_csa_tree_lt_140_15_groupi_n_20, lbl5_en1_csa_tree_lt_140_15_groupi_n_21, lbl5_en1_csa_tree_lt_140_15_groupi_n_22, lbl5_en1_csa_tree_lt_140_15_groupi_n_23 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_24, lbl5_en1_csa_tree_lt_140_15_groupi_n_25, lbl5_en1_csa_tree_lt_140_15_groupi_n_26, lbl5_en1_csa_tree_lt_140_15_groupi_n_27, lbl5_en1_csa_tree_lt_140_15_groupi_n_28 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_29, lbl5_en1_csa_tree_lt_140_15_groupi_n_30, lbl5_en1_csa_tree_lt_140_15_groupi_n_31, lbl5_en1_csa_tree_lt_140_15_groupi_n_32, lbl5_en1_csa_tree_lt_140_15_groupi_n_33 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_34, lbl5_en1_csa_tree_lt_140_15_groupi_n_36, lbl5_en1_csa_tree_lt_140_15_groupi_n_37, lbl5_en1_csa_tree_lt_140_15_groupi_n_38, lbl5_en1_csa_tree_lt_140_15_groupi_n_39 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_40, lbl5_en1_csa_tree_lt_140_15_groupi_n_41, lbl5_en1_csa_tree_lt_140_15_groupi_n_42, lbl5_en1_csa_tree_lt_140_15_groupi_n_43, lbl5_en1_csa_tree_lt_140_15_groupi_n_44 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_45, lbl5_en1_csa_tree_lt_140_15_groupi_n_46, lbl5_en1_csa_tree_lt_140_15_groupi_n_47, lbl5_en1_csa_tree_lt_140_15_groupi_n_48, lbl5_en1_csa_tree_lt_140_15_groupi_n_49 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_50, lbl5_en1_csa_tree_lt_140_15_groupi_n_51, lbl5_en1_csa_tree_lt_140_15_groupi_n_52, lbl5_en1_csa_tree_lt_140_15_groupi_n_53, lbl5_en1_csa_tree_lt_140_15_groupi_n_54 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_55, lbl5_en1_csa_tree_lt_140_15_groupi_n_56, lbl5_en1_csa_tree_lt_140_15_groupi_n_57, lbl5_en1_csa_tree_lt_140_15_groupi_n_58, lbl5_en1_csa_tree_lt_140_15_groupi_n_59 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_60, lbl5_en1_csa_tree_lt_140_15_groupi_n_61, lbl5_en1_csa_tree_lt_140_15_groupi_n_62, lbl5_en1_csa_tree_lt_140_15_groupi_n_63, lbl5_en1_csa_tree_lt_140_15_groupi_n_64 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_65, lbl5_en1_csa_tree_lt_140_15_groupi_n_66, lbl5_en1_csa_tree_lt_140_15_groupi_n_67, lbl5_en1_csa_tree_lt_140_15_groupi_n_68, lbl5_en1_csa_tree_lt_140_15_groupi_n_69 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_112, lbl5_en1_csa_tree_lt_140_15_groupi_n_114, lbl5_en1_csa_tree_lt_140_15_groupi_n_118, lbl5_en1_csa_tree_lt_140_15_groupi_n_119, lbl5_en1_csa_tree_lt_140_15_groupi_n_120 : std_logic;
  signal lbl5_en1_csa_tree_lt_140_15_groupi_n_121, lbl5_en1_csa_tree_lt_140_15_groupi_n_123, lbl5_en1_csa_tree_lt_140_15_groupi_n_124, lbl5_en1_frozen_boost, lbl5_en1_inc_add_127_23_n_0 : std_logic;
  signal lbl5_en1_inc_add_127_23_n_2, lbl5_en1_inc_add_127_23_n_4, lbl5_en1_inc_add_127_23_n_6, lbl5_en1_inc_add_127_23_n_8, lbl5_en1_inc_add_127_23_n_10 : std_logic;
  signal lbl5_en1_inc_add_127_23_n_12, lbl5_en1_inc_add_127_23_n_14, lbl5_en1_inc_add_127_23_n_16, lbl5_en1_inc_add_127_23_n_18, lbl5_en1_inc_add_127_23_n_20 : std_logic;
  signal lbl5_en1_inc_add_127_23_n_22, lbl5_en1_inc_add_127_23_n_24, lbl5_en1_inc_add_127_23_n_26, lbl5_en1_inc_add_127_23_n_28, lbl5_en1_inc_add_127_23_n_30 : std_logic;
  signal lbl5_en1_inc_add_127_23_n_32, lbl5_en1_n_0, lbl5_en1_n_1, lbl5_en1_n_2, lbl5_en1_n_3 : std_logic;
  signal lbl5_en1_n_4, lbl5_en1_n_5, lbl5_en1_n_6, lbl5_en1_n_7, lbl5_en1_n_8 : std_logic;
  signal lbl5_en1_n_9, lbl5_en1_n_10, lbl5_en1_n_11, lbl5_en1_n_12, lbl5_en1_n_13 : std_logic;
  signal lbl5_en1_n_14, lbl5_en1_n_15, lbl5_en1_n_16, lbl5_en1_n_17, lbl5_en1_n_18 : std_logic;
  signal lbl5_en1_n_19, lbl5_en1_n_20, lbl5_en1_n_21, lbl5_en1_n_22, lbl5_en1_n_23 : std_logic;
  signal lbl5_en1_n_24, lbl5_en1_n_25, lbl5_en1_n_26, lbl5_en1_n_27, lbl5_en1_n_28 : std_logic;
  signal lbl5_en1_n_29, lbl5_en1_n_30, lbl5_en1_n_31, lbl5_en1_n_32, lbl5_en1_n_33 : std_logic;
  signal lbl5_en1_n_34, lbl5_en1_n_35, lbl5_en1_n_36, lbl5_en1_n_37, lbl5_en1_n_38 : std_logic;
  signal lbl5_en1_n_39, lbl5_en1_n_40, lbl5_en1_n_41, lbl5_en1_n_42, lbl5_en1_n_43 : std_logic;
  signal lbl5_en1_n_44, lbl5_en1_n_45, lbl5_en1_n_46, lbl5_en1_n_47, lbl5_en1_n_48 : std_logic;
  signal lbl5_en1_n_49, lbl5_en1_n_50, lbl5_en1_n_51, lbl5_en1_n_52, lbl5_en1_n_53 : std_logic;
  signal lbl5_en1_n_54, lbl5_en1_n_55, lbl5_en1_n_56, lbl5_en1_n_57, lbl5_en1_n_58 : std_logic;
  signal lbl5_en1_n_59, lbl5_en1_n_60, lbl5_en1_n_61, lbl5_en1_n_62, lbl5_en1_n_63 : std_logic;
  signal lbl5_en1_n_64, lbl5_en1_n_65, lbl5_en1_n_66, lbl5_en1_n_67, lbl5_en1_n_68 : std_logic;
  signal lbl5_en1_n_69, lbl5_en1_n_70, lbl5_en1_n_71, lbl5_en1_n_72, lbl5_en1_n_73 : std_logic;
  signal lbl5_en1_n_74, lbl5_en1_n_75, lbl5_en1_n_76, lbl5_en1_n_77, lbl5_en1_n_78 : std_logic;
  signal lbl5_en1_n_79, lbl5_en1_n_80, lbl5_en1_n_81, lbl5_en1_n_82, lbl5_en1_n_83 : std_logic;
  signal lbl5_en1_n_84, lbl5_en1_n_85, lbl5_en1_n_86, lbl5_en1_n_87, lbl5_en1_n_88 : std_logic;
  signal lbl5_en1_n_89, lbl5_en1_n_90, lbl5_en1_n_91, lbl5_en1_n_92, lbl5_en1_n_93 : std_logic;
  signal lbl5_en1_n_94, lbl5_en1_n_95, lbl5_en1_n_96, lbl5_en1_n_97, lbl5_en1_n_98 : std_logic;
  signal lbl5_en1_n_99, lbl5_en1_n_100, lbl5_en1_n_101, lbl5_en1_n_102, lbl5_en1_n_103 : std_logic;
  signal lbl5_en1_n_104, lbl5_en1_n_105, lbl5_en1_n_106, lbl5_en1_n_107, lbl5_en1_n_108 : std_logic;
  signal lbl5_en1_n_109, lbl5_en1_n_110, lbl5_en1_n_111, lbl5_en1_n_112, lbl5_en1_n_113 : std_logic;
  signal lbl5_en1_n_114, lbl5_en1_n_115, lbl5_en1_n_116, lbl5_en1_n_117, lbl5_en1_n_118 : std_logic;
  signal lbl5_en1_n_119, lbl5_en1_n_120, lbl5_en1_n_121, lbl5_en1_n_122, lbl5_en1_n_123 : std_logic;
  signal lbl5_en1_n_124, lbl5_en1_n_125, lbl5_en1_n_126, lbl5_en1_n_127, lbl5_en1_n_128 : std_logic;
  signal lbl5_en1_n_129, lbl5_en1_n_130, lbl5_en1_n_131, lbl5_en1_n_132, lbl5_en1_n_133 : std_logic;
  signal lbl5_en1_n_134, lbl5_en1_n_135, lbl5_en1_n_136, lbl5_en1_n_137, lbl5_en1_n_138 : std_logic;
  signal lbl5_en1_n_139, lbl5_en1_n_140, lbl5_en1_n_141, lbl5_en1_n_142, lbl5_en1_n_143 : std_logic;
  signal lbl5_en1_n_144, lbl5_en1_n_145, lbl5_en1_n_146, lbl5_en1_n_147, lbl5_en1_n_148 : std_logic;
  signal lbl5_en1_n_149, lbl5_en1_n_150, lbl5_en1_n_151, lbl5_en1_n_152, lbl5_en1_n_153 : std_logic;
  signal lbl5_en1_n_154, lbl5_en1_n_155, lbl5_en1_n_156, lbl5_en1_n_157, lbl5_en1_n_158 : std_logic;
  signal lbl5_en1_n_159, lbl5_en1_n_160, lbl5_en1_n_161, lbl5_en1_n_162, lbl5_en1_n_163 : std_logic;
  signal lbl5_en1_n_164, lbl5_en1_n_165, lbl5_en1_n_166, lbl5_en1_n_167, lbl5_en1_n_168 : std_logic;
  signal lbl5_en1_n_169, lbl5_en1_n_170, lbl5_en1_n_171, lbl5_en1_n_172, lbl5_en1_n_173 : std_logic;
  signal lbl5_en1_n_174, lbl5_en1_n_175, lbl5_en1_n_176, lbl5_en1_n_177, lbl5_en1_n_178 : std_logic;
  signal lbl5_en1_n_179, lbl5_en1_n_180, lbl5_en1_n_181, lbl5_en1_n_182, lbl5_en1_n_183 : std_logic;
  signal lbl5_en1_n_186, lbl5_en1_n_190, lbl5_en1_n_191, lbl5_en1_n_192, lbl5_en1_n_194 : std_logic;
  signal lbl5_en1_n_195, lbl5_en1_n_197, lbl5_en1_n_200, lbl5_en1_n_202, lbl5_en1_n_203 : std_logic;
  signal lbl5_en1_n_204, lbl5_en1_n_205, lbl5_en1_n_206, lbl5_en1_n_207, lbl5_en1_n_208 : std_logic;
  signal lbl5_en1_n_209, lbl5_en1_n_210, lbl5_en1_n_211, lbl5_en1_n_212, lbl5_en1_n_213 : std_logic;
  signal lbl5_en1_n_214, lbl5_en1_n_215, lbl5_en1_n_216, lbl5_en1_n_217, lbl5_en1_n_218 : std_logic;
  signal lbl5_en1_n_219, lbl5_en1_n_220, lbl5_en1_n_222, lbl5_en1_n_223, lbl5_en1_n_224 : std_logic;
  signal lbl5_en1_n_225, lbl5_en1_n_226, lbl5_en1_n_227, lbl5_en1_n_228, lbl5_en1_n_229 : std_logic;
  signal lbl5_en1_n_230, lbl5_en1_n_231, lbl5_en1_n_232, lbl5_en1_n_233, lbl5_en1_n_234 : std_logic;
  signal lbl5_en1_n_235, lbl5_en1_n_236, lbl5_en1_n_237, lbl5_en1_n_238, lbl5_en1_n_239 : std_logic;
  signal lbl5_en1_n_240, lbl5_en1_n_241, lbl5_en1_n_242, lbl5_en1_n_243, lbl5_en1_n_244 : std_logic;
  signal lbl5_en1_n_245, lbl5_en1_n_246, lbl5_en1_n_247, lbl5_en1_n_248, lbl5_en1_n_249 : std_logic;
  signal lbl5_en1_n_250, lbl5_en1_n_251, lbl5_en1_n_252, lbl5_en1_n_253, lbl5_en1_n_254 : std_logic;
  signal lbl5_en1_n_255, lbl5_en1_n_256, lbl5_en1_n_257, lbl5_en1_n_258, lbl5_en1_n_259 : std_logic;
  signal lbl5_en1_n_260, lbl5_en1_n_261, lbl5_en1_n_262, lbl5_en1_n_263, lbl5_en1_n_264 : std_logic;
  signal lbl5_en1_n_265, lbl5_en1_n_267, lbl5_en1_n_268, lbl5_en1_n_269, lbl5_en1_n_270 : std_logic;
  signal lbl5_en1_n_271, lbl5_en1_n_272, lbl5_en1_n_273, lbl5_en1_n_274, lbl5_en1_n_275 : std_logic;
  signal lbl5_en1_n_276, lbl5_en1_n_277, lbl5_en1_n_278, lbl5_en1_n_280, lbl5_en1_n_281 : std_logic;
  signal lbl5_en1_n_282, lbl5_en1_n_284, lbl5_en1_n_285, lbl5_en1_n_286, lbl5_en1_n_287 : std_logic;
  signal lbl5_en1_n_288, lbl5_en1_n_289, lbl5_en1_n_290, lbl5_en1_n_291, lbl5_en1_n_292 : std_logic;
  signal lbl5_en1_n_293, lbl5_en1_n_294, lbl5_en1_n_295, lbl5_en1_n_296, lbl5_en1_n_297 : std_logic;
  signal lbl5_en1_n_298, lbl5_en1_n_299, lbl5_en1_n_300, lbl5_en1_n_301, lbl5_en1_n_302 : std_logic;
  signal lbl5_en1_n_303, lbl5_en1_n_304, lbl5_en1_n_305, lbl5_en1_n_306, lbl5_en1_n_307 : std_logic;
  signal lbl5_en1_n_308, lbl5_en1_n_309, lbl5_en1_n_310, lbl5_en1_n_311, lbl5_en1_n_312 : std_logic;
  signal lbl5_en1_n_313, lbl5_en1_n_314, lbl5_en1_n_315, lbl5_en1_n_316, lbl5_en1_n_317 : std_logic;
  signal lbl5_en1_n_318, lbl5_en1_n_319, lbl5_en1_n_320, lbl5_en1_n_331, lbl5_en1_n_332 : std_logic;
  signal lbl5_en1_n_333, lbl5_en1_prev_crash, lbl5_en1_prev_engine, lbl5_engine_en, lbl5_expl_n_1 : std_logic;
  signal lbl5_n_0, lbl5_n_2, memory_ready, pulse_audio, reset_vga_mem : std_logic;
  signal start_between, write_enable, x_increment, y_increment : std_logic;

begin

  FE_PHC349_lbl5_en1_new_period_17 : DEL01BWP7T port map(I => FE_PHN349_lbl5_en1_new_period_17, Z => FE_PHN322_lbl5_en1_new_period_17);
  FE_PHC348_lbl5_en1_new_period_1 : CKBD0BWP7T port map(I => lbl5_en1_new_period(1), Z => FE_PHN348_lbl5_en1_new_period_1);
  FE_PHC347_lbl5_en1_new_period_3 : DEL01BWP7T port map(I => FE_PHN319_lbl5_en1_new_period_3, Z => FE_PHN347_lbl5_en1_new_period_3);
  FE_PHC346_lbl5_en1_n_10 : DEL01BWP7T port map(I => FE_PHN320_lbl5_en1_n_10, Z => FE_PHN346_lbl5_en1_n_10);
  FE_PHC345_lbl5_en1_new_period_5 : DEL01BWP7T port map(I => FE_PHN250_lbl5_en1_new_period_5, Z => FE_PHN345_lbl5_en1_new_period_5);
  FE_PHC344_lbl5_en1_n_301 : DEL01BWP7T port map(I => lbl5_en1_n_301, Z => FE_PHN344_lbl5_en1_n_301);
  FE_PHC343_lbl1_cm_n_8 : DEL01BWP7T port map(I => FE_PHN343_lbl1_cm_n_8, Z => lbl1_cm_n_8);
  FE_PHC342_lbl1_rw_n_84 : DEL01BWP7T port map(I => lbl1_rw_n_84, Z => FE_PHN342_lbl1_rw_n_84);
  FE_PHC341_lbl5_en0_new_period_6 : DEL0BWP7T port map(I => FE_PHN341_lbl5_en0_new_period_6, Z => lbl5_en0_new_period(6));
  FE_PHC340_lbl0_border_1 : DEL01BWP7T port map(I => FE_PHN155_lbl0_border_1, Z => FE_PHN340_lbl0_border_1);
  FE_PHC339_lbl1_cm_state_0 : DEL01BWP7T port map(I => lbl1_cm_state(0), Z => FE_PHN339_lbl1_cm_state_0);
  FE_PHC338_lbl5_en0_period_7 : DEL01BWP7T port map(I => FE_PHN145_lbl5_en0_period_7, Z => FE_PHN338_lbl5_en0_period_7);
  FE_PHC337_lbl5_en1_new_period_0 : DEL0BWP7T port map(I => lbl5_en1_new_period(0), Z => FE_PHN337_lbl5_en1_new_period_0);
  FE_PHC336_lbl2_v_count_7 : DEL01BWP7T port map(I => FE_PHN194_lbl2_v_count_7, Z => FE_PHN336_lbl2_v_count_7);
  FE_PHC335_lbl1_cur_w_1 : DEL01BWP7T port map(I => lbl1_cur_w(1), Z => FE_PHN335_lbl1_cur_w_1);
  FE_PHC334_lbl5_en1_new_period_4 : DEL0BWP7T port map(I => lbl5_en1_new_period(4), Z => FE_PHN334_lbl5_en1_new_period_4);
  FE_PHC333_lbl0_mem_com_state_2 : DEL01BWP7T port map(I => lbl0_mem_com_state(2), Z => FE_PHN333_lbl0_mem_com_state_2);
  FE_PHC332_lbl1_cur_w_3 : DEL01BWP7T port map(I => FE_PHN332_lbl1_cur_w_3, Z => FE_PHN208_lbl1_cur_w_3);
  FE_PHC331_lbl5_en1_new_period_5 : CKBD0BWP7T port map(I => lbl5_en1_new_period(5), Z => FE_PHN331_lbl5_en1_new_period_5);
  FE_PHC330_lbl0_border_0 : DEL01BWP7T port map(I => lbl0_border_0, Z => FE_PHN330_lbl0_border_0);
  FE_PHC329_lbl5_en0_n_7 : DEL01BWP7T port map(I => FE_PHN329_lbl5_en0_n_7, Z => FE_PHN232_lbl5_en0_n_7);
  FE_PHC328_direction_in_2 : DEL01BWP7T port map(I => FE_PHN151_direction_in_2, Z => FE_PHN328_direction_in_2);
  FE_PHC327_lbl5_en1_n_3 : DEL01BWP7T port map(I => lbl5_en1_n_3, Z => FE_PHN327_lbl5_en1_n_3);
  FE_PHC326_lbl1_cur_w_5 : DEL01BWP7T port map(I => FE_PHN326_lbl1_cur_w_5, Z => FE_PHN187_lbl1_cur_w_5);
  FE_PHC325_lbl5_en1_count_6 : DEL01BWP7T port map(I => lbl5_en1_count(6), Z => FE_PHN325_lbl5_en1_count_6);
  FE_PHC324_y_address_0 : DEL01BWP7T port map(I => y_address(0), Z => FE_PHN324_y_address_0);
  FE_PHC323_lbl2_jumps_synced_7 : DEL01BWP7T port map(I => FE_PHN143_lbl2_jumps_synced_7, Z => FE_PHN323_lbl2_jumps_synced_7);
  FE_PHC322_lbl5_en1_new_period_17 : CKBD0BWP7T port map(I => FE_PHN322_lbl5_en1_new_period_17, Z => FE_PHN136_lbl5_en1_new_period_17);
  FE_PHC321_lbl5_en1_new_period_1 : DEL02BWP7T port map(I => FE_PHN348_lbl5_en1_new_period_1, Z => FE_PHN321_lbl5_en1_new_period_1);
  FE_PHC320_lbl5_en1_n_10 : CKBD0BWP7T port map(I => FE_PHN245_lbl5_en1_n_10, Z => FE_PHN320_lbl5_en1_n_10);
  FE_PHC319_lbl5_en1_new_period_3 : CKBD0BWP7T port map(I => lbl5_en1_new_period(3), Z => FE_PHN319_lbl5_en1_new_period_3);
  FE_PHC318_lbl5_en0_new_period_5 : DEL0BWP7T port map(I => FE_PHN249_lbl5_en0_new_period_5, Z => FE_PHN318_lbl5_en0_new_period_5);
  FE_PHC317_lbl5_en1_new_period_14 : CKBD0BWP7T port map(I => FE_PHN221_lbl5_en1_new_period_14, Z => FE_PHN317_lbl5_en1_new_period_14);
  FE_PHC316_lbl2_v_count_9 : CKBD0BWP7T port map(I => FE_PHN238_lbl2_v_count_9, Z => FE_PHN316_lbl2_v_count_9);
  FE_PHC315_lbl0_busy_count_0 : DEL0BWP7T port map(I => FE_PHN258_lbl0_busy_count_0, Z => FE_PHN315_lbl0_busy_count_0);
  FE_PHC314_lbl0_mem_com_state_0 : CKBD0BWP7T port map(I => lbl0_mem_com_state(0), Z => FE_PHN314_lbl0_mem_com_state_0);
  FE_PHC313_lbl5_en1_frozen_bits_1 : DEL01BWP7T port map(I => lbl5_en1_frozen_bits(1), Z => FE_PHN313_lbl5_en1_frozen_bits_1);
  FE_PHC312_lbl5_en1_new_period_8 : CKBD0BWP7T port map(I => FE_PHN216_lbl5_en1_new_period_8, Z => FE_PHN312_lbl5_en1_new_period_8);
  FE_PHC311_lbl0_n_47 : DEL0BWP7T port map(I => lbl0_n_47, Z => FE_PHN311_lbl0_n_47);
  FE_PHC310_lbl1_cy_n_10 : BUFFD2BWP7T port map(I => lbl1_cy_n_10, Z => FE_PHN310_lbl1_cy_n_10);
  FE_PHC309_lbl0_n_539 : DEL01BWP7T port map(I => lbl0_n_539, Z => FE_PHN309_lbl0_n_539);
  FE_PHC308_lbl1_cm_n_23 : CKBD0BWP7T port map(I => lbl1_cm_n_23, Z => FE_PHN308_lbl1_cm_n_23);
  FE_PHC307_lbl0_n_46 : CKBD0BWP7T port map(I => lbl0_n_46, Z => FE_PHN307_lbl0_n_46);
  FE_PHC306_lbl5_en1_n_178 : CKBD0BWP7T port map(I => FE_PHN306_lbl5_en1_n_178, Z => lbl5_en1_n_178);
  FE_PHC305_lbl1_cy_n_3 : CKBD0BWP7T port map(I => lbl1_cy_n_3, Z => FE_PHN305_lbl1_cy_n_3);
  FE_PHC304_lbl1_cex_n_3 : DEL0BWP7T port map(I => lbl1_cex_n_3, Z => FE_PHN304_lbl1_cex_n_3);
  FE_PHC303_lbl1_cey_n_3 : DEL0BWP7T port map(I => FE_PHN303_lbl1_cey_n_3, Z => lbl1_cey_n_3);
  FE_PHC302_lbl1_cy_n_7 : DEL01BWP7T port map(I => lbl1_cy_n_7, Z => FE_PHN302_lbl1_cy_n_7);
  FE_PHC301_lbl1_cy_n_5 : DEL01BWP7T port map(I => lbl1_cy_n_5, Z => FE_PHN301_lbl1_cy_n_5);
  FE_PHC300_lbl1_cx_n_10 : DEL0BWP7T port map(I => lbl1_cx_n_10, Z => FE_PHN300_lbl1_cx_n_10);
  FE_PHC299_lbl1_cw_n_7 : DEL1BWP7T port map(I => lbl1_cw_n_7, Z => FE_PHN299_lbl1_cw_n_7);
  FE_PHC298_lbl1_cx_n_7 : DEL01BWP7T port map(I => lbl1_cx_n_7, Z => FE_PHN298_lbl1_cx_n_7);
  FE_PHC297_lbl1_cw_n_16 : DEL1BWP7T port map(I => lbl1_cw_n_16, Z => FE_PHN297_lbl1_cw_n_16);
  FE_PHC296_lbl1_cx_n_5 : DEL01BWP7T port map(I => lbl1_cx_n_5, Z => FE_PHN296_lbl1_cx_n_5);
  FE_PHC295_lbl5_expl_n_1 : DEL0BWP7T port map(I => lbl5_expl_n_1, Z => FE_PHN295_lbl5_expl_n_1);
  FE_PHC294_lbl0_n_34 : DEL0BWP7T port map(I => lbl0_n_34, Z => FE_PHN294_lbl0_n_34);
  FE_PHC293_lbl1_cm_n_24 : DEL0BWP7T port map(I => lbl1_cm_n_24, Z => FE_PHN293_lbl1_cm_n_24);
  FE_PHC292_lbl5_en0_n_46 : DEL0BWP7T port map(I => lbl5_en0_n_46, Z => FE_PHN292_lbl5_en0_n_46);
  FE_PHC291_lbl1_rw_n_68 : CKBD0BWP7T port map(I => lbl1_rw_n_68, Z => FE_PHN291_lbl1_rw_n_68);
  FE_PHC290_lbl5_en1_n_300 : DEL0BWP7T port map(I => lbl5_en1_n_300, Z => FE_PHN290_lbl5_en1_n_300);
  FE_PHC289_lbl5_en1_n_179 : DEL0BWP7T port map(I => lbl5_en1_n_179, Z => FE_PHN289_lbl5_en1_n_179);
  FE_PHC288_lbl1_cw_n_3 : DEL0BWP7T port map(I => lbl1_cw_n_3, Z => FE_PHN288_lbl1_cw_n_3);
  FE_PHC287_lbl5_en1_n_183 : DEL0BWP7T port map(I => lbl5_en1_n_183, Z => FE_PHN287_lbl5_en1_n_183);
  FE_PHC286_lbl5_en0_n_296 : DEL0BWP7T port map(I => FE_PHN286_lbl5_en0_n_296, Z => lbl5_en0_n_296);
  FE_PHC285_lbl5_en0_n_157 : DEL1BWP7T port map(I => FE_PHN285_lbl5_en0_n_157, Z => lbl5_en0_n_157);
  FE_PHC284_lbl5_en0_n_156 : DEL0BWP7T port map(I => lbl5_en0_n_156, Z => FE_PHN284_lbl5_en0_n_156);
  FE_PHC283_lbl1_cx_n_3 : CKBD0BWP7T port map(I => lbl1_cx_n_3, Z => FE_PHN283_lbl1_cx_n_3);
  FE_PHC282_lbl5_en0_n_161 : DEL0BWP7T port map(I => FE_PHN282_lbl5_en0_n_161, Z => lbl5_en0_n_161);
  FE_PHC281_lbl5_en0_n_298 : DEL0BWP7T port map(I => lbl5_en0_n_298, Z => FE_PHN281_lbl5_en0_n_298);
  FE_PHC280_lbl5_en1_n_302 : DEL0BWP7T port map(I => FE_PHN280_lbl5_en1_n_302, Z => lbl5_en1_n_302);
  FE_PHC279_lbl0_n_37 : DEL1BWP7T port map(I => lbl0_n_37, Z => FE_PHN279_lbl0_n_37);
  FE_PHC278_lbl5_en1_n_182 : DEL1BWP7T port map(I => FE_PHN278_lbl5_en1_n_182, Z => lbl5_en1_n_182);
  FE_PHC277_lbl1_cey_n_1 : DEL1BWP7T port map(I => lbl1_cey_n_1, Z => FE_PHN277_lbl1_cey_n_1);
  FE_PHC276_lbl0_n_43 : DEL0BWP7T port map(I => lbl0_n_43, Z => FE_PHN276_lbl0_n_43);
  FE_PHC275_lbl1_cex_n_1 : DEL1BWP7T port map(I => lbl1_cex_n_1, Z => FE_PHN275_lbl1_cex_n_1);
  FE_PHC274_lbl0_n_38 : DEL0BWP7T port map(I => lbl0_n_38, Z => FE_PHN274_lbl0_n_38);
  FE_PHC273_lbl5_en1_n_280 : DEL0BWP7T port map(I => lbl5_en1_n_280, Z => FE_PHN273_lbl5_en1_n_280);
  FE_PHC272_lbl0_n_42 : DEL0BWP7T port map(I => lbl0_n_42, Z => FE_PHN272_lbl0_n_42);
  FE_PHC271_lbl5_en0_n_276 : DEL0BWP7T port map(I => lbl5_en0_n_276, Z => FE_PHN271_lbl5_en0_n_276);
  FE_PHC270_lbl5_en0_n_155 : DEL0BWP7T port map(I => lbl5_en0_n_155, Z => FE_PHN270_lbl5_en0_n_155);
  FE_PHC269_lbl0_n_45 : DEL1BWP7T port map(I => lbl0_n_45, Z => FE_PHN269_lbl0_n_45);
  FE_PHC268_lbl0_n_44 : DEL1BWP7T port map(I => lbl0_n_44, Z => FE_PHN268_lbl0_n_44);
  FE_PHC267_lbl5_en0_n_158 : DEL1BWP7T port map(I => FE_PHN267_lbl5_en0_n_158, Z => lbl5_en0_n_158);
  FE_PHC266_lbl0_mem_com_state_0 : DEL02BWP7T port map(I => FE_PHN266_lbl0_mem_com_state_0, Z => lbl0_mem_com_state(0));
  FE_PHC265_lbl5_en0_new_period_6 : DEL1BWP7T port map(I => lbl5_en0_new_period(6), Z => FE_PHN265_lbl5_en0_new_period_6);
  FE_PHC264_lbl5_en0_period_18 : DEL0BWP7T port map(I => FE_PHN264_lbl5_en0_period_18, Z => lbl5_en0_period(18));
  FE_PHC263_lbl5_en0_period_16 : DEL0BWP7T port map(I => lbl5_en0_period(16), Z => FE_PHN263_lbl5_en0_period_16);
  FE_PHC262_lbl0_mem_com_state_3 : CKBD0BWP7T port map(I => lbl0_mem_com_state(3), Z => FE_PHN262_lbl0_mem_com_state_3);
  FE_PHC261_lbl5_en0_period_17 : DEL1BWP7T port map(I => FE_PHN261_lbl5_en0_period_17, Z => lbl5_en0_period(17));
  FE_PHC260_lbl5_en1_period_17 : DEL1BWP7T port map(I => FE_PHN260_lbl5_en1_period_17, Z => lbl5_en1_period(17));
  FE_PHC259_lbl5_en1_period_16 : DEL0BWP7T port map(I => lbl5_en1_period(16), Z => FE_PHN259_lbl5_en1_period_16);
  FE_PHC258_lbl0_busy_count_0 : DEL02BWP7T port map(I => lbl0_busy_count(0), Z => FE_PHN258_lbl0_busy_count_0);
  FE_PHC257_x_address_3 : DEL02BWP7T port map(I => FE_PHN257_x_address_3, Z => x_address(3));
  FE_PHC256_lbl0_mem_com_state_1 : CKBD0BWP7T port map(I => FE_PHN256_lbl0_mem_com_state_1, Z => lbl0_mem_com_state(1));
  FE_PHC255_direction_0_1 : DEL1BWP7T port map(I => direction_0(1), Z => FE_PHN255_direction_0_1);
  FE_PHC254_lbl5_en0_count_16 : DEL02BWP7T port map(I => FE_PHN254_lbl5_en0_count_16, Z => lbl5_en0_count(16));
  FE_PHC253_direction_between_3 : DEL01BWP7T port map(I => direction_between(3), Z => FE_PHN253_direction_between_3);
  FE_PHC252_lbl5_en1_new_period_1 : DEL02BWP7T port map(I => FE_PHN252_lbl5_en1_new_period_1, Z => lbl5_en1_new_period(1));
  FE_PHC251_lbl5_en0_count_17 : DEL1BWP7T port map(I => FE_PHN251_lbl5_en0_count_17, Z => lbl5_en0_count(17));
  FE_PHC250_lbl5_en1_new_period_5 : DEL02BWP7T port map(I => FE_PHN331_lbl5_en1_new_period_5, Z => FE_PHN250_lbl5_en1_new_period_5);
  FE_PHC249_lbl5_en0_new_period_5 : DEL02BWP7T port map(I => lbl5_en0_new_period(5), Z => FE_PHN249_lbl5_en0_new_period_5);
  FE_PHC248_lbl5_en1_new_period_3 : DEL02BWP7T port map(I => FE_PHN248_lbl5_en1_new_period_3, Z => lbl5_en1_new_period(3));
  FE_PHC247_y_address_3 : CKBD0BWP7T port map(I => y_address(3), Z => FE_PHN247_y_address_3);
  FE_PHC246_lbl5_en0_new_period_2 : DEL1BWP7T port map(I => FE_PHN246_lbl5_en0_new_period_2, Z => lbl5_en0_new_period(2));
  FE_PHC245_lbl5_en1_n_10 : DEL02BWP7T port map(I => lbl5_en1_n_10, Z => FE_PHN245_lbl5_en1_n_10);
  FE_PHC244_lbl5_en1_new_period_2 : DEL1BWP7T port map(I => lbl5_en1_new_period(2), Z => FE_PHN244_lbl5_en1_new_period_2);
  FE_PHC243_lbl5_en0_new_period_14 : DEL0BWP7T port map(I => FE_PHN243_lbl5_en0_new_period_14, Z => lbl5_en0_new_period(14));
  FE_PHC242_lbl5_en0_new_period_4 : DEL1BWP7T port map(I => FE_PHN242_lbl5_en0_new_period_4, Z => lbl5_en0_new_period(4));
  FE_PHC241_direction_between_2 : DEL01BWP7T port map(I => direction_between(2), Z => FE_PHN241_direction_between_2);
  FE_PHC240_direction_between_0 : CKBD0BWP7T port map(I => direction_between(0), Z => FE_PHN240_direction_between_0);
  FE_PHC239_lbl5_en1_new_period_7 : DEL02BWP7T port map(I => lbl5_en1_new_period(7), Z => FE_PHN239_lbl5_en1_new_period_7);
  FE_PHC238_lbl2_v_count_9 : DEL02BWP7T port map(I => lbl2_v_count(9), Z => FE_PHN238_lbl2_v_count_9);
  FE_PHC237_lbl5_en0_new_period_8 : DEL0BWP7T port map(I => lbl5_en0_new_period(8), Z => FE_PHN237_lbl5_en0_new_period_8);
  FE_PHC236_lbl5_en0_new_period_13 : DEL0BWP7T port map(I => lbl5_en0_new_period(13), Z => FE_PHN236_lbl5_en0_new_period_13);
  FE_PHC235_read_memory_in_4 : CKBD0BWP7T port map(I => read_memory_in(4), Z => FE_PHN235_read_memory_in_4);
  FE_PHC234_lbl5_en0_new_period_10 : DEL0BWP7T port map(I => lbl5_en0_new_period(10), Z => FE_PHN234_lbl5_en0_new_period_10);
  FE_PHC233_lbl5_en0_new_period_11 : DEL1BWP7T port map(I => lbl5_en0_new_period(11), Z => FE_PHN233_lbl5_en0_new_period_11);
  FE_PHC232_lbl5_en0_n_7 : DEL02BWP7T port map(I => FE_PHN232_lbl5_en0_n_7, Z => lbl5_en0_n_7);
  FE_PHC231_read_memory_in_5 : CKBD0BWP7T port map(I => read_memory_in(5), Z => FE_PHN231_read_memory_in_5);
  FE_PHC230_lbl5_en0_new_period_9 : DEL1BWP7T port map(I => FE_PHN230_lbl5_en0_new_period_9, Z => lbl5_en0_new_period(9));
  FE_PHC229_lbl2_n_21 : DEL01BWP7T port map(I => lbl2_n_21, Z => FE_PHN229_lbl2_n_21);
  FE_PHC228_lbl5_en1_new_period_13 : DEL1BWP7T port map(I => lbl5_en1_new_period(13), Z => FE_PHN228_lbl5_en1_new_period_13);
  FE_PHC227_lbl5_en1_n_4 : DEL1BWP7T port map(I => lbl5_en1_n_4, Z => FE_PHN227_lbl5_en1_n_4);
  FE_PHC226_lbl5_en1_n_2 : DEL1BWP7T port map(I => lbl5_en1_n_2, Z => FE_PHN226_lbl5_en1_n_2);
  FE_PHC225_lbl5_en1_new_period_4 : DEL02BWP7T port map(I => FE_PHN334_lbl5_en1_new_period_4, Z => FE_PHN225_lbl5_en1_new_period_4);
  FE_PHC224_lbl5_en1_n_3 : DEL02BWP7T port map(I => FE_PHN327_lbl5_en1_n_3, Z => FE_PHN224_lbl5_en1_n_3);
  FE_PHC223_lbl5_en1_n_8 : DEL0BWP7T port map(I => lbl5_en1_n_8, Z => FE_PHN223_lbl5_en1_n_8);
  FE_PHC222_lbl5_en1_n_9 : DEL01BWP7T port map(I => lbl5_en1_n_9, Z => FE_PHN222_lbl5_en1_n_9);
  FE_PHC221_lbl5_en1_new_period_14 : DEL02BWP7T port map(I => lbl5_en1_new_period(14), Z => FE_PHN221_lbl5_en1_new_period_14);
  FE_PHC220_lbl5_en0_new_period_7 : DEL0BWP7T port map(I => FE_PHN220_lbl5_en0_new_period_7, Z => lbl5_en0_new_period(7));
  FE_PHC219_lbl5_en0_new_period_0 : DEL1BWP7T port map(I => FE_PHN219_lbl5_en0_new_period_0, Z => lbl5_en0_new_period(0));
  FE_PHC218_direction_between_1 : DEL01BWP7T port map(I => direction_between(1), Z => FE_PHN218_direction_between_1);
  FE_PHC217_read_memory_in_0 : BUFFD2BWP7T port map(I => read_memory_in(0), Z => FE_PHN217_read_memory_in_0);
  FE_PHC216_lbl5_en1_new_period_8 : DEL02BWP7T port map(I => lbl5_en1_new_period(8), Z => FE_PHN216_lbl5_en1_new_period_8);
  FE_PHC215_lbl5_en1_new_period_9 : DEL2BWP7T port map(I => FE_PHN215_lbl5_en1_new_period_9, Z => lbl5_en1_new_period(9));
  FE_PHC214_lbl1_cur_w_1 : DEL02BWP7T port map(I => FE_PHN335_lbl1_cur_w_1, Z => FE_PHN214_lbl1_cur_w_1);
  FE_PHC213_lbl5_en1_new_period_16 : DEL0BWP7T port map(I => lbl5_en1_new_period(16), Z => FE_PHN213_lbl5_en1_new_period_16);
  FE_PHC212_lbl1_cur_w_2 : DEL02BWP7T port map(I => lbl1_cur_w(2), Z => FE_PHN212_lbl1_cur_w_2);
  FE_PHC211_lbl5_en1_new_period_0 : DEL02BWP7T port map(I => FE_PHN337_lbl5_en1_new_period_0, Z => FE_PHN211_lbl5_en1_new_period_0);
  FE_PHC210_lbl0_n_65 : DEL01BWP7T port map(I => lbl0_n_65, Z => FE_PHN210_lbl0_n_65);
  FE_PHC209_lbl5_en1_n_6 : DEL0BWP7T port map(I => FE_PHN209_lbl5_en1_n_6, Z => lbl5_en1_n_6);
  FE_PHC208_lbl1_cur_w_3 : DEL02BWP7T port map(I => FE_PHN208_lbl1_cur_w_3, Z => lbl1_cur_w(3));
  FE_PHC207_lbl0_n_81 : DEL01BWP7T port map(I => lbl0_n_81, Z => FE_PHN207_lbl0_n_81);
  FE_PHC206_lbl5_en1_new_period_11 : DEL1BWP7T port map(I => lbl5_en1_new_period(11), Z => FE_PHN206_lbl5_en1_new_period_11);
  FE_PHC205_read_memory_in_1 : CKBD0BWP7T port map(I => read_memory_in(1), Z => FE_PHN205_read_memory_in_1);
  FE_PHC204_lbl5_en1_n_7 : DEL0BWP7T port map(I => FE_PHN204_lbl5_en1_n_7, Z => lbl5_en1_n_7);
  FE_PHC203_lbl5_en1_new_period_15 : DEL0BWP7T port map(I => lbl5_en1_new_period(15), Z => FE_PHN203_lbl5_en1_new_period_15);
  FE_PHC202_lbl5_en0_new_period_15 : DEL0BWP7T port map(I => FE_PHN202_lbl5_en0_new_period_15, Z => lbl5_en0_new_period(15));
  FE_PHC201_read_memory_in_2 : CKBD0BWP7T port map(I => read_memory_in(2), Z => FE_PHN201_read_memory_in_2);
  FE_PHC200_lbl1_cur_w_0 : DEL0BWP7T port map(I => lbl1_cur_w(0), Z => FE_PHN200_lbl1_cur_w_0);
  FE_PHC199_lbl5_en0_frozen_boost : DEL01BWP7T port map(I => lbl5_en0_frozen_boost, Z => FE_PHN199_lbl5_en0_frozen_boost);
  FE_PHC198_read_memory_in_6 : CKBD0BWP7T port map(I => read_memory_in(6), Z => FE_PHN198_read_memory_in_6);
  FE_PHC197_lbl1_cur_w_4 : DEL0BWP7T port map(I => FE_PHN197_lbl1_cur_w_4, Z => lbl1_cur_w(4));
  FE_PHC196_lbl0_next_direction_0_1 : DEL01BWP7T port map(I => lbl0_next_direction_0(1), Z => FE_PHN196_lbl0_next_direction_0_1);
  FE_PHC195_lbl5_en1_n_290 : CKBD0BWP7T port map(I => lbl5_en1_n_290, Z => FE_PHN195_lbl5_en1_n_290);
  FE_PHC194_lbl2_v_count_7 : CKBD0BWP7T port map(I => lbl2_v_count(7), Z => FE_PHN194_lbl2_v_count_7);
  FE_PHC193_read_memory_in_7 : CKBD0BWP7T port map(I => read_memory_in(7), Z => FE_PHN193_read_memory_in_7);
  FE_PHC192_lbl5_en0_new_period_16 : DEL0BWP7T port map(I => FE_PHN192_lbl5_en0_new_period_16, Z => lbl5_en0_new_period(16));
  FE_PHC191_lbl1_cur_w_6 : DEL0BWP7T port map(I => FE_PHN191_lbl1_cur_w_6, Z => lbl1_cur_w(6));
  FE_PHC190_lbl5_en1_n_285 : DEL0BWP7T port map(I => FE_PHN190_lbl5_en1_n_285, Z => lbl5_en1_n_285);
  FE_PHC189_lbl5_en1_n_292 : CKBD4BWP7T port map(I => lbl5_en1_n_292, Z => FE_PHN189_lbl5_en1_n_292);
  FE_PHC188_lbl5_en0_n_281 : DEL0BWP7T port map(I => lbl5_en0_n_281, Z => FE_PHN188_lbl5_en0_n_281);
  FE_PHC187_lbl1_cur_w_5 : DEL02BWP7T port map(I => FE_PHN187_lbl1_cur_w_5, Z => lbl1_cur_w(5));
  FE_PHC186_lbl1_rw_n_0 : DEL01BWP7T port map(I => lbl1_rw_n_0, Z => FE_PHN186_lbl1_rw_n_0);
  FE_PHC185_lbl5_en1_count_17 : DEL02BWP7T port map(I => lbl5_en1_count(17), Z => FE_PHN185_lbl5_en1_count_17);
  FE_PHC184_lbl5_en0_n_285 : DEL0BWP7T port map(I => lbl5_en0_n_285, Z => FE_PHN184_lbl5_en0_n_285);
  FE_PHC183_lbl5_en1_n_288 : DEL0BWP7T port map(I => lbl5_en1_n_288, Z => FE_PHN183_lbl5_en1_n_288);
  FE_PHC182_lbl0_counter_busy_counter_state_0 : DEL0BWP7T port map(I => lbl0_counter_busy_counter_state(0), Z => FE_PHN182_lbl0_counter_busy_counter_state_0);
  FE_PHC181_lbl5_en0_n_283 : DEL0BWP7T port map(I => FE_PHN181_lbl5_en0_n_283, Z => lbl5_en0_n_283);
  FE_PHC180_lbl5_en0_n_289 : DEL0BWP7T port map(I => lbl5_en0_n_289, Z => FE_PHN180_lbl5_en0_n_289);
  FE_PHC179_lbl5_en1_n_287 : DEL0BWP7T port map(I => lbl5_en1_n_287, Z => FE_PHN179_lbl5_en1_n_287);
  FE_PHC178_lbl5_en1_n_289 : DEL0BWP7T port map(I => lbl5_en1_n_289, Z => FE_PHN178_lbl5_en1_n_289);
  FE_PHC177_lbl5_en0_n_282 : DEL0BWP7T port map(I => lbl5_en0_n_282, Z => FE_PHN177_lbl5_en0_n_282);
  FE_PHC176_lbl5_en0_n_290 : DEL0BWP7T port map(I => lbl5_en0_n_290, Z => FE_PHN176_lbl5_en0_n_290);
  FE_PHC175_lbl5_en0_n_291 : DEL0BWP7T port map(I => lbl5_en0_n_291, Z => FE_PHN175_lbl5_en0_n_291);
  FE_PHC174_lbl1_cm_n_52 : DEL0BWP7T port map(I => FE_PHN174_lbl1_cm_n_52, Z => lbl1_cm_n_52);
  FE_PHC173_lbl5_en1_n_293 : CKBD3BWP7T port map(I => lbl5_en1_n_293, Z => FE_PHN173_lbl5_en1_n_293);
  FE_PHC172_lbl5_en0_n_293 : DEL0BWP7T port map(I => FE_PHN172_lbl5_en0_n_293, Z => lbl5_en0_n_293);
  FE_PHC171_direction_0_0 : DEL1BWP7T port map(I => direction_0(0), Z => FE_PHN171_direction_0_0);
  FE_PHC170_lbl5_en1_n_295 : DEL0BWP7T port map(I => FE_PHN170_lbl5_en1_n_295, Z => lbl5_en1_n_295);
  FE_PHC169_lbl5_en0_n_288 : BUFFD3BWP7T port map(I => lbl5_en0_n_288, Z => FE_PHN169_lbl5_en0_n_288);
  FE_PHC168_lbl5_en0_n_287 : DEL0BWP7T port map(I => FE_PHN168_lbl5_en0_n_287, Z => lbl5_en0_n_287);
  FE_PHC167_lbl0_n_63 : DEL01BWP7T port map(I => lbl0_n_63, Z => FE_PHN167_lbl0_n_63);
  FE_PHC166_lbl5_en0_n_286 : BUFFD3BWP7T port map(I => lbl5_en0_n_286, Z => FE_PHN166_lbl5_en0_n_286);
  FE_PHC165_lbl5_en0_n_284 : BUFFD3BWP7T port map(I => lbl5_en0_n_284, Z => FE_PHN165_lbl5_en0_n_284);
  FE_PHC164_lbl0_counter_busy_counter_state_1 : DEL1BWP7T port map(I => FE_PHN164_lbl0_counter_busy_counter_state_1, Z => lbl0_counter_busy_counter_state(1));
  FE_PHC163_lbl0_border_0 : CKBD0BWP7T port map(I => FE_PHN330_lbl0_border_0, Z => FE_PHN163_lbl0_border_0);
  FE_PHC162_lbl5_en1_n_298 : DEL0BWP7T port map(I => lbl5_en1_n_298, Z => FE_PHN162_lbl5_en1_n_298);
  FE_PHC161_lbl5_en1_n_294 : DEL0BWP7T port map(I => lbl5_en1_n_294, Z => FE_PHN161_lbl5_en1_n_294);
  FE_PHC160_lbl5_en0_n_292 : DEL0BWP7T port map(I => FE_PHN160_lbl5_en0_n_292, Z => lbl5_en0_n_292);
  FE_PHC159_lbl5_en1_n_291 : DEL0BWP7T port map(I => lbl5_en1_n_291, Z => FE_PHN159_lbl5_en1_n_291);
  FE_PHC158_lbl5_en0_n_294 : DEL0BWP7T port map(I => lbl5_en0_n_294, Z => FE_PHN158_lbl5_en0_n_294);
  FE_PHC157_lbl1_cex_n_4 : DEL0BWP7T port map(I => lbl1_cex_n_4, Z => FE_PHN157_lbl1_cex_n_4);
  FE_PHC156_lbl1_cm_n_22 : DEL0BWP7T port map(I => FE_PHN156_lbl1_cm_n_22, Z => lbl1_cm_n_22);
  FE_PHC155_lbl0_border_1 : CKBD0BWP7T port map(I => lbl0_border_1, Z => FE_PHN155_lbl0_border_1);
  FE_PHC154_lbl1_cey_n_4 : DEL0BWP7T port map(I => lbl1_cey_n_4, Z => FE_PHN154_lbl1_cey_n_4);
  FE_PHC153_read_memory_in_3 : CKBD0BWP7T port map(I => read_memory_in(3), Z => FE_PHN153_read_memory_in_3);
  FE_PHC152_lbl1_rw_n_27 : DEL01BWP7T port map(I => lbl1_rw_n_27, Z => FE_PHN152_lbl1_rw_n_27);
  FE_PHC151_direction_in_2 : DEL0BWP7T port map(I => direction_in(2), Z => FE_PHN151_direction_in_2);
  FE_PHC150_lbl2_v_count_8 : CKBD0BWP7T port map(I => lbl2_v_count(8), Z => FE_PHN150_lbl2_v_count_8);
  FE_PHC149_lbl1_rw_n_58 : DEL0BWP7T port map(I => lbl1_rw_n_58, Z => FE_PHN149_lbl1_rw_n_58);
  FE_PHC148_lbl5_en1_n_296 : DEL0BWP7T port map(I => lbl5_en1_n_296, Z => FE_PHN148_lbl5_en1_n_296);
  FE_PHC147_lbl5_en1_period_4 : DEL0BWP7T port map(I => lbl5_en1_period(4), Z => FE_PHN147_lbl5_en1_period_4);
  FE_PHC146_lbl5_en1_n_5 : DEL1BWP7T port map(I => lbl5_en1_n_5, Z => FE_PHN146_lbl5_en1_n_5);
  FE_PHC145_lbl5_en0_period_7 : DEL0BWP7T port map(I => lbl5_en0_period(7), Z => FE_PHN145_lbl5_en0_period_7);
  FE_PHC144_lbl5_en0_period_13 : DEL0BWP7T port map(I => lbl5_en0_period(13), Z => FE_PHN144_lbl5_en0_period_13);
  FE_PHC143_lbl2_jumps_synced_7 : DEL0BWP7T port map(I => lbl2_jumps_synced(7), Z => FE_PHN143_lbl2_jumps_synced_7);
  FE_PHC142_boost_audio_1 : DEL0BWP7T port map(I => boost_audio_1, Z => FE_PHN142_boost_audio_1);
  FE_PHC141_lbl5_en0_n_295 : DEL0BWP7T port map(I => lbl5_en0_n_295, Z => FE_PHN141_lbl5_en0_n_295);
  FE_PHC140_lbl5_en1_frozen_boost : CKBD0BWP7T port map(I => lbl5_en1_frozen_boost, Z => FE_PHN140_lbl5_en1_frozen_boost);
  FE_PHC139_lbl5_en1_n_299 : DEL0BWP7T port map(I => FE_PHN139_lbl5_en1_n_299, Z => lbl5_en1_n_299);
  FE_PHC138_lbl2_v_count_6 : CKBD0BWP7T port map(I => lbl2_v_count(6), Z => FE_PHN138_lbl2_v_count_6);
  FE_PHC137_lbl5_en1_count_16 : DEL02BWP7T port map(I => lbl5_en1_count(16), Z => FE_PHN137_lbl5_en1_count_16);
  FE_PHC136_lbl5_en1_new_period_17 : DEL02BWP7T port map(I => FE_PHN136_lbl5_en1_new_period_17, Z => lbl5_en1_new_period(17));
  FE_PHC135_lbl5_en1_n_297 : DEL0BWP7T port map(I => lbl5_en1_n_297, Z => FE_PHN135_lbl5_en1_n_297);
  FE_PHC134_direction_in_0 : DEL1BWP7T port map(I => direction_in(0), Z => FE_PHN134_direction_in_0);
  FE_PHC133_lbl2_data_synced_2 : DEL0BWP7T port map(I => lbl2_data_synced(2), Z => FE_PHN133_lbl2_data_synced_2);
  FE_PHC132_lbl5_en0_period_10 : DEL1BWP7T port map(I => lbl5_en0_period(10), Z => FE_PHN132_lbl5_en0_period_10);
  FE_PHC131_lbl5_en1_frozen_bits_0 : DEL1BWP7T port map(I => lbl5_en1_frozen_bits(0), Z => FE_PHN131_lbl5_en1_frozen_bits_0);
  FE_PHC130_lbl5_en1_n_286 : CKBD0BWP7T port map(I => lbl5_en1_n_286, Z => FE_PHN130_lbl5_en1_n_286);
  FE_PHC129_lbl2_data_synced_1 : DEL0BWP7T port map(I => lbl2_data_synced(1), Z => FE_PHN129_lbl2_data_synced_1);
  FE_PHC128_direction_1_1 : DEL1BWP7T port map(I => direction_1(1), Z => FE_PHN128_direction_1_1);
  FE_PHC127_direction_in_1 : DEL1BWP7T port map(I => direction_in(1), Z => FE_PHN127_direction_in_1);
  FE_PHC126_direction_1_0 : DEL1BWP7T port map(I => direction_1(0), Z => FE_PHN126_direction_1_0);
  FE_PHC125_lbl5_en1_frozen_bits_1 : DEL0BWP7T port map(I => FE_PHN125_lbl5_en1_frozen_bits_1, Z => lbl5_en1_frozen_bits(1));
  FE_PHC124_lbl5_en0_period_5 : DEL0BWP7T port map(I => lbl5_en0_period(5), Z => FE_PHN124_lbl5_en0_period_5);
  FE_PHC123_lbl5_en1_period_6 : DEL1BWP7T port map(I => lbl5_en1_period(6), Z => FE_PHN123_lbl5_en1_period_6);
  FE_PHC122_lbl2_data_synced_5 : DEL0BWP7T port map(I => lbl2_data_synced(5), Z => FE_PHN122_lbl2_data_synced_5);
  FE_PHC121_lbl5_en0_frozen_bits_2 : DEL1BWP7T port map(I => FE_PHN121_lbl5_en0_frozen_bits_2, Z => lbl5_en0_frozen_bits(2));
  FE_PHC120_lbl2_data_synced_6 : DEL0BWP7T port map(I => lbl2_data_synced(6), Z => FE_PHN120_lbl2_data_synced_6);
  FE_PHC119_lbl5_en1_period_5 : DEL1BWP7T port map(I => lbl5_en1_period(5), Z => FE_PHN119_lbl5_en1_period_5);
  FE_PHC118_lbl5_en0_n_6 : DEL0BWP7T port map(I => lbl5_en0_n_6, Z => FE_PHN118_lbl5_en0_n_6);
  FE_PHC117_lbl5_en1_n_13 : DEL1BWP7T port map(I => lbl5_en1_n_13, Z => FE_PHN117_lbl5_en1_n_13);
  FE_PHC116_lbl2_data_synced_0 : DEL0BWP7T port map(I => lbl2_data_synced(0), Z => FE_PHN116_lbl2_data_synced_0);
  FE_PHC115_lbl5_en0_period_9 : DEL1BWP7T port map(I => lbl5_en0_period(9), Z => FE_PHN115_lbl5_en0_period_9);
  FE_PHC114_lbl5_en1_period_9 : DEL1BWP7T port map(I => lbl5_en1_period(9), Z => FE_PHN114_lbl5_en1_period_9);
  FE_PHC113_lbl5_en1_period_7 : DEL1BWP7T port map(I => lbl5_en1_period(7), Z => FE_PHN113_lbl5_en1_period_7);
  FE_PHC112_lbl5_en1_period_12 : DEL1BWP7T port map(I => lbl5_en1_period(12), Z => FE_PHN112_lbl5_en1_period_12);
  FE_PHC111_lbl5_en0_n_8 : DEL0BWP7T port map(I => lbl5_en0_n_8, Z => FE_PHN111_lbl5_en0_n_8);
  FE_PHC110_lbl5_en0_period_3 : DEL1BWP7T port map(I => lbl5_en0_period(3), Z => FE_PHN110_lbl5_en0_period_3);
  FE_PHC109_lbl2_data_synced_4 : DEL0BWP7T port map(I => lbl2_data_synced(4), Z => FE_PHN109_lbl2_data_synced_4);
  FE_PHC108_lbl5_en0_frozen_bits_3 : DEL1BWP7T port map(I => FE_PHN108_lbl5_en0_frozen_bits_3, Z => lbl5_en0_frozen_bits(3));
  FE_PHC107_lbl5_en0_period_14 : DEL0BWP7T port map(I => lbl5_en0_period(14), Z => FE_PHN107_lbl5_en0_period_14);
  FE_PHC106_lbl5_en1_period_10 : DEL1BWP7T port map(I => lbl5_en1_period(10), Z => FE_PHN106_lbl5_en1_period_10);
  FE_PHC105_lbl5_en0_period_12 : DEL1BWP7T port map(I => lbl5_en0_period(12), Z => FE_PHN105_lbl5_en0_period_12);
  FE_PHC104_boost_audio_0 : DEL0BWP7T port map(I => boost_audio_0, Z => FE_PHN104_boost_audio_0);
  FE_PHC103_direction_in_3 : DEL1BWP7T port map(I => direction_in(3), Z => FE_PHN103_direction_in_3);
  FE_PHC102_lbl5_en1_period_11 : DEL1BWP7T port map(I => lbl5_en1_period(11), Z => FE_PHN102_lbl5_en1_period_11);
  FE_PHC101_lbl2_data_synced_3 : DEL0BWP7T port map(I => lbl2_data_synced(3), Z => FE_PHN101_lbl2_data_synced_3);
  FE_PHC100_lbl5_en0_n_5 : DEL0BWP7T port map(I => lbl5_en0_n_5, Z => FE_PHN100_lbl5_en0_n_5);
  FE_PHC99_lbl5_en1_period_1 : DEL0BWP7T port map(I => lbl5_en1_period(1), Z => FE_PHN99_lbl5_en1_period_1);
  FE_PHC98_lbl5_en0_period_2 : DEL0BWP7T port map(I => lbl5_en0_period(2), Z => FE_PHN98_lbl5_en0_period_2);
  FE_PHC97_lbl5_en0_period_8 : DEL0BWP7T port map(I => lbl5_en0_period(8), Z => FE_PHN97_lbl5_en0_period_8);
  FE_PHC96_lbl5_en1_frozen_bits_3 : DEL1BWP7T port map(I => FE_PHN96_lbl5_en1_frozen_bits_3, Z => lbl5_en1_frozen_bits(3));
  FE_PHC95_lbl5_en1_period_13 : DEL0BWP7T port map(I => lbl5_en1_period(13), Z => FE_PHN95_lbl5_en1_period_13);
  FE_PHC94_lbl2_borders_synced_1 : DEL1BWP7T port map(I => lbl2_borders_synced(1), Z => FE_PHN94_lbl2_borders_synced_1);
  FE_PHC93_lbl2_borders_synced_5 : DEL1BWP7T port map(I => lbl2_borders_synced(5), Z => FE_PHN93_lbl2_borders_synced_5);
  FE_PHC92_lbl5_en0_period_6 : DEL0BWP7T port map(I => lbl5_en0_period(6), Z => FE_PHN92_lbl5_en0_period_6);
  FE_PHC91_lbl5_en0_period_15 : DEL0BWP7T port map(I => lbl5_en0_period(15), Z => FE_PHN91_lbl5_en0_period_15);
  FE_PHC90_lbl5_en1_period_14 : DEL0BWP7T port map(I => lbl5_en1_period(14), Z => FE_PHN90_lbl5_en1_period_14);
  FE_PHC89_lbl5_en1_period_8 : DEL0BWP7T port map(I => lbl5_en1_period(8), Z => FE_PHN89_lbl5_en1_period_8);
  FE_PHC88_lbl5_en0_period_0 : DEL0BWP7T port map(I => lbl5_en0_period(0), Z => FE_PHN88_lbl5_en0_period_0);
  FE_PHC87_lbl5_en1_period_18 : DEL0BWP7T port map(I => lbl5_en1_period(18), Z => FE_PHN87_lbl5_en1_period_18);
  FE_PHC86_lbl5_en1_period_0 : DEL0BWP7T port map(I => lbl5_en1_period(0), Z => FE_PHN86_lbl5_en1_period_0);
  FE_PHC85_lbl2_borders_synced_6 : DEL1BWP7T port map(I => lbl2_borders_synced(6), Z => FE_PHN85_lbl2_borders_synced_6);
  FE_PHC84_lbl5_en1_period_15 : DEL0BWP7T port map(I => lbl5_en1_period(15), Z => FE_PHN84_lbl5_en1_period_15);
  FE_PHC83_lbl2_borders_synced_2 : DEL1BWP7T port map(I => lbl2_borders_synced(2), Z => FE_PHN83_lbl2_borders_synced_2);
  FE_PHC82_lbl2_borders_synced_7 : DEL1BWP7T port map(I => lbl2_borders_synced(7), Z => FE_PHN82_lbl2_borders_synced_7);
  FE_PHC81_lbl5_en1_frozen_bits_2 : DEL1BWP7T port map(I => lbl5_en1_frozen_bits(2), Z => FE_PHN81_lbl5_en1_frozen_bits_2);
  FE_PHC80_lbl5_en0_period_4 : DEL0BWP7T port map(I => lbl5_en0_period(4), Z => FE_PHN80_lbl5_en0_period_4);
  FE_PHC79_lbl2_data_synced_7 : DEL0BWP7T port map(I => lbl2_data_synced(7), Z => FE_PHN79_lbl2_data_synced_7);
  FE_PHC78_lbl2_jumps_synced_5 : DEL1BWP7T port map(I => lbl2_jumps_synced(5), Z => FE_PHN78_lbl2_jumps_synced_5);
  FE_PHC77_lbl2_jumps_synced_3 : DEL1BWP7T port map(I => lbl2_jumps_synced(3), Z => FE_PHN77_lbl2_jumps_synced_3);
  FE_PHC76_lbl2_jumps_synced_6 : DEL1BWP7T port map(I => lbl2_jumps_synced(6), Z => FE_PHN76_lbl2_jumps_synced_6);
  FE_PHC75_lbl2_jumps_synced_0 : DEL1BWP7T port map(I => lbl2_jumps_synced(0), Z => FE_PHN75_lbl2_jumps_synced_0);
  FE_PHC74_lbl2_borders_synced_4 : DEL1BWP7T port map(I => lbl2_borders_synced(4), Z => FE_PHN74_lbl2_borders_synced_4);
  FE_PHC73_lbl2_borders_synced_3 : DEL1BWP7T port map(I => lbl2_borders_synced(3), Z => FE_PHN73_lbl2_borders_synced_3);
  FE_PHC72_lbl5_en0_period_11 : DEL0BWP7T port map(I => lbl5_en0_period(11), Z => FE_PHN72_lbl5_en0_period_11);
  FE_PHC71_lbl2_jumps_synced_1 : DEL1BWP7T port map(I => lbl2_jumps_synced(1), Z => FE_PHN71_lbl2_jumps_synced_1);
  FE_PHC70_lbl5_en1_period_2 : DEL0BWP7T port map(I => lbl5_en1_period(2), Z => FE_PHN70_lbl5_en1_period_2);
  FE_PHC69_lbl2_jumps_synced_4 : DEL1BWP7T port map(I => lbl2_jumps_synced(4), Z => FE_PHN69_lbl2_jumps_synced_4);
  FE_PHC68_lbl2_borders_synced_0 : DEL1BWP7T port map(I => lbl2_borders_synced(0), Z => FE_PHN68_lbl2_borders_synced_0);
  FE_PHC67_lbl2_jumps_synced_2 : DEL1BWP7T port map(I => lbl2_jumps_synced(2), Z => FE_PHN67_lbl2_jumps_synced_2);
  FE_PHC66_lbl5_en1_period_3 : DEL0BWP7T port map(I => lbl5_en1_period(3), Z => FE_PHN66_lbl5_en1_period_3);
  FE_PHC65_start_in : DEL0BWP7T port map(I => start_in, Z => FE_PHN65_start_in);
  FE_PHC64_lbl5_en0_new_period_17 : DEL2BWP7T port map(I => lbl5_en0_new_period(17), Z => FE_PHN64_lbl5_en0_new_period_17);
  FE_PHC63_lbl5_en0_period_1 : DEL0BWP7T port map(I => lbl5_en0_period(1), Z => FE_PHN63_lbl5_en0_period_1);
  FE_PHC62_lbl5_en0_n_12 : DEL0BWP7T port map(I => lbl5_en0_n_12, Z => FE_PHN62_lbl5_en0_n_12);
  FE_PHC61_lbl0_booster_sync : DEL0BWP7T port map(I => lbl0_booster_sync, Z => FE_PHN61_lbl0_booster_sync);
  FE_PHC60_lbl5_expl_shifter_15 : DEL1BWP7T port map(I => FE_PHN60_lbl5_expl_shifter_15, Z => lbl5_expl_shifter(15));
  FE_PHC59_lbl5_expl_shifter_21 : DEL1BWP7T port map(I => lbl5_expl_shifter(21), Z => FE_PHN59_lbl5_expl_shifter_21);
  FE_PHC58_lbl5_expl_shifter_6 : DEL1BWP7T port map(I => FE_PHN58_lbl5_expl_shifter_6, Z => lbl5_expl_shifter(6));
  FE_PHC57_lbl5_en0_frozen_bits_0 : DEL1BWP7T port map(I => FE_PHN57_lbl5_en0_frozen_bits_0, Z => lbl5_en0_frozen_bits(0));
  FE_PHC56_lbl5_en0_n_16 : CKBD0BWP7T port map(I => lbl5_en0_n_16, Z => FE_PHN56_lbl5_en0_n_16);
  FE_PHC55_lbl3_temp1_1 : DEL2BWP7T port map(I => lbl3_temp1(1), Z => FE_PHN55_lbl3_temp1_1);
  FE_PHC54_lbl5_en0_n_11 : DEL1BWP7T port map(I => FE_PHN54_lbl5_en0_n_11, Z => lbl5_en0_n_11);
  FE_PHC53_lbl5_en0_frozen_bits_1 : DEL1BWP7T port map(I => lbl5_en0_frozen_bits(1), Z => FE_PHN53_lbl5_en0_frozen_bits_1);
  FE_PHC52_lbl5_en0_n_14 : DEL0BWP7T port map(I => lbl5_en0_n_14, Z => FE_PHN52_lbl5_en0_n_14);
  FE_PHC51_lbl5_en0_n_9 : DEL0BWP7T port map(I => lbl5_en0_n_9, Z => FE_PHN51_lbl5_en0_n_9);
  FE_PHC50_lbl3_temp2 : DEL1BWP7T port map(I => lbl3_temp2, Z => FE_PHN50_lbl3_temp2);
  FE_PHC49_lbl5_expl_shifter_20 : DEL1BWP7T port map(I => lbl5_expl_shifter(20), Z => FE_PHN49_lbl5_expl_shifter_20);
  FE_PHC48_lbl3_temp1_0 : DEL1BWP7T port map(I => lbl3_temp1(0), Z => FE_PHN48_lbl3_temp1_0);
  FE_PHC47_lbl5_expl_shifter_4 : DEL1BWP7T port map(I => lbl5_expl_shifter(4), Z => FE_PHN47_lbl5_expl_shifter_4);
  FE_PHC46_lbl5_expl_shifter_22 : DEL1BWP7T port map(I => lbl5_expl_shifter(22), Z => FE_PHN46_lbl5_expl_shifter_22);
  FE_PHC45_lbl5_expl_shifter_17 : DEL1BWP7T port map(I => lbl5_expl_shifter(17), Z => FE_PHN45_lbl5_expl_shifter_17);
  FE_PHC44_lbl5_expl_shifter_16 : DEL1BWP7T port map(I => lbl5_expl_shifter(16), Z => FE_PHN44_lbl5_expl_shifter_16);
  FE_PHC43_lbl5_expl_shifter_7 : DEL1BWP7T port map(I => FE_PHN43_lbl5_expl_shifter_7, Z => lbl5_expl_shifter(7));
  FE_PHC42_lbl5_expl_shifter_5 : DEL1BWP7T port map(I => FE_PHN42_lbl5_expl_shifter_5, Z => lbl5_expl_shifter(5));
  FE_PHC41_lbl5_expl_shifter_13 : DEL1BWP7T port map(I => lbl5_expl_shifter(13), Z => FE_PHN41_lbl5_expl_shifter_13);
  FE_PHC40_lbl5_expl_shifter_11 : DEL1BWP7T port map(I => FE_PHN40_lbl5_expl_shifter_11, Z => lbl5_expl_shifter(11));
  FE_PHC39_lbl5_expl_shifter_14 : DEL1BWP7T port map(I => lbl5_expl_shifter(14), Z => FE_PHN39_lbl5_expl_shifter_14);
  FE_PHC38_lbl5_expl_shifter_10 : DEL1BWP7T port map(I => FE_PHN38_lbl5_expl_shifter_10, Z => lbl5_expl_shifter(10));
  FE_PHC37_lbl5_expl_shifter_12 : DEL1BWP7T port map(I => FE_PHN37_lbl5_expl_shifter_12, Z => lbl5_expl_shifter(12));
  FE_PHC36_lbl5_expl_shifter_9 : DEL1BWP7T port map(I => lbl5_expl_shifter(9), Z => FE_PHN36_lbl5_expl_shifter_9);
  FE_PHC35_lbl5_expl_shifter_8 : DEL1BWP7T port map(I => lbl5_expl_shifter(8), Z => FE_PHN35_lbl5_expl_shifter_8);
  FE_PHC34_lbl5_expl_shifter_18 : DEL1BWP7T port map(I => FE_PHN34_lbl5_expl_shifter_18, Z => lbl5_expl_shifter(18));
  FE_PHC33_lbl5_expl_shifter_19 : DEL1BWP7T port map(I => lbl5_expl_shifter(19), Z => FE_PHN33_lbl5_expl_shifter_19);
  FE_PHC32_lbl3_temp1_3 : DEL1BWP7T port map(I => FE_PHN32_lbl3_temp1_3, Z => lbl3_temp1(3));
  FE_PHC31_lbl5_en1_new_period_18 : DEL1BWP7T port map(I => FE_PHN31_lbl5_en1_new_period_18, Z => lbl5_en1_new_period(18));
  FE_PHC30_lbl5_en0_new_period_18 : DEL1BWP7T port map(I => FE_PHN30_lbl5_en0_new_period_18, Z => lbl5_en0_new_period(18));
  FE_PHC29_lbl3_temp1_2 : DEL1BWP7T port map(I => FE_PHN29_lbl3_temp1_2, Z => lbl3_temp1(2));
  FE_PHC28_lbl5_bits_3 : DEL1BWP7T port map(I => FE_PHN28_lbl5_bits_3, Z => lbl5_bits(3));
  FE_PHC27_lbl5_bits_2 : DEL1BWP7T port map(I => FE_PHN27_lbl5_bits_2, Z => lbl5_bits(2));
  FE_PHC26_lbl5_bits_0 : DEL1BWP7T port map(I => lbl5_bits(0), Z => FE_PHN26_lbl5_bits_0);
  FE_PHC25_lbl5_bits_1 : DEL1BWP7T port map(I => lbl5_bits(1), Z => FE_PHN25_lbl5_bits_1);
  FE_OFC5_FE_DBTN24_rst : BUFFD2BWP7T port map(I => FE_DBTN24_rst, Z => FE_OFN5_FE_DBTN24_rst);
  FE_OFC4_memory_enable_out : BUFFD5BWP7T port map(I => FE_OFN4_memory_enable_out, Z => memory_enable_out);
  FE_OFC1_rst : DEL01BWP7T port map(I => rst, Z => FE_OFN1_rst);
  FE_OFC0_lbl2_n_2 : CKBD1BWP7T port map(I => lbl2_n_2, Z => FE_OFN0_lbl2_n_2);
  CTS_ccl_a_BUF_clk_G0_L2_4 : CKBD10BWP7T port map(I => CTS_22, Z => CTS_21);
  CTS_ccl_a_BUF_clk_G0_L2_3 : CKBD10BWP7T port map(I => CTS_22, Z => CTS_20);
  CTS_ccl_a_BUF_clk_G0_L2_2 : CKBD10BWP7T port map(I => CTS_22, Z => CTS_19);
  CTS_ccl_a_BUF_clk_G0_L2_1 : CKBD10BWP7T port map(I => CTS_22, Z => CTS_18);
  CTS_ccl_a_BUF_clk_G0_L1_1 : CKBD10BWP7T port map(I => clk, Z => CTS_22);
  FE_DBTC24_rst : CKND1BWP7T port map(I => FE_OFN1_rst, ZN => FE_DBTN24_rst);
  FE_DBTC23_memory_reset_out : INVD1BWP7T port map(I => memory_reset_out, ZN => FE_DBTN23_memory_reset_out);
  FE_DBTC22_position_1_10 : INVD1BWP7T port map(I => position_1(10), ZN => FE_DBTN22_position_1_10);
  FE_DBTC21_lbl2_h_count_3 : INVD1BWP7T port map(I => lbl2_h_count(3), ZN => FE_DBTN21_lbl2_h_count_3);
  FE_DBTC20_lbl2_h_count_2 : INVD0BWP7T port map(I => lbl2_h_count(2), ZN => FE_DBTN20_lbl2_h_count_2);
  FE_DBTC19_lbl2_h_count_1 : INVD0BWP7T port map(I => lbl2_h_count(1), ZN => FE_DBTN19_lbl2_h_count_1);
  FE_DBTC18_lbl2_v_count_2 : INVD1BWP7T port map(I => lbl2_v_count(2), ZN => FE_DBTN18_lbl2_v_count_2);
  FE_DBTC17_lbl5_en0_n_301 : INVD0BWP7T port map(I => lbl5_en0_n_301, ZN => FE_DBTN17_lbl5_en0_n_301);
  FE_DBTC16_lbl5_en0_n_304 : INVD1BWP7T port map(I => lbl5_en0_n_304, ZN => FE_DBTN16_lbl5_en0_n_304);
  FE_DBTC15_lbl5_en0_n_306 : INVD1BWP7T port map(I => lbl5_en0_n_306, ZN => FE_DBTN15_lbl5_en0_n_306);
  FE_DBTC14_lbl5_en0_n_305 : INVD1BWP7T port map(I => lbl5_en0_n_305, ZN => FE_DBTN14_lbl5_en0_n_305);
  FE_DBTC13_lbl5_en0_n_309 : INVD1BWP7T port map(I => lbl5_en0_n_309, ZN => FE_DBTN13_lbl5_en0_n_309);
  FE_DBTC12_lbl5_en0_n_303 : INVD1BWP7T port map(I => lbl5_en0_n_303, ZN => FE_DBTN12_lbl5_en0_n_303);
  FE_DBTC11_lbl5_en0_n_308 : INVD1BWP7T port map(I => lbl5_en0_n_308, ZN => FE_DBTN11_lbl5_en0_n_308);
  FE_DBTC10_lbl5_en0_n_311 : INVD1BWP7T port map(I => lbl5_en0_n_311, ZN => FE_DBTN10_lbl5_en0_n_311);
  FE_DBTC9_lbl5_en0_n_302 : INVD1BWP7T port map(I => lbl5_en0_n_302, ZN => FE_DBTN9_lbl5_en0_n_302);
  FE_DBTC8_lbl5_en1_n_305 : INVD0BWP7T port map(I => lbl5_en1_n_305, ZN => FE_DBTN8_lbl5_en1_n_305);
  FE_DBTC7_lbl5_en1_n_308 : INVD1BWP7T port map(I => lbl5_en1_n_308, ZN => FE_DBTN7_lbl5_en1_n_308);
  FE_DBTC6_lbl5_en1_n_310 : INVD1BWP7T port map(I => lbl5_en1_n_310, ZN => FE_DBTN6_lbl5_en1_n_310);
  FE_DBTC5_lbl5_en1_n_309 : INVD1BWP7T port map(I => lbl5_en1_n_309, ZN => FE_DBTN5_lbl5_en1_n_309);
  FE_DBTC4_lbl5_en1_n_313 : INVD1BWP7T port map(I => lbl5_en1_n_313, ZN => FE_DBTN4_lbl5_en1_n_313);
  FE_DBTC3_lbl5_en1_n_307 : INVD1BWP7T port map(I => lbl5_en1_n_307, ZN => FE_DBTN3_lbl5_en1_n_307);
  FE_DBTC2_lbl5_en1_n_312 : INVD1BWP7T port map(I => lbl5_en1_n_312, ZN => FE_DBTN2_lbl5_en1_n_312);
  FE_DBTC1_lbl5_en1_n_315 : INVD1BWP7T port map(I => lbl5_en1_n_315, ZN => FE_DBTN1_lbl5_en1_n_315);
  FE_DBTC0_lbl5_en1_n_306 : INVD1BWP7T port map(I => lbl5_en1_n_306, ZN => FE_DBTN0_lbl5_en1_n_306);
  lbl2_g2832 : NR4D0BWP7T port map(A1 => lbl2_n_142, A2 => lbl2_n_53, A3 => lbl2_n_124, A4 => lbl2_n_113, ZN => lbl2_n_190);
  lbl2_g2833 : NR4D0BWP7T port map(A1 => lbl2_n_141, A2 => lbl2_n_53, A3 => lbl2_n_125, A4 => lbl2_n_114, ZN => lbl2_n_189);
  lbl2_g2834 : ND4D0BWP7T port map(A1 => lbl2_n_140, A2 => lbl2_n_127, A3 => lbl2_n_120, A4 => lbl2_n_117, ZN => lbl2_n_142);
  lbl2_g2835 : ND4D0BWP7T port map(A1 => lbl2_n_139, A2 => lbl2_n_130, A3 => lbl2_n_118, A4 => lbl2_n_119, ZN => lbl2_n_141);
  lbl2_g2836 : NR3D0BWP7T port map(A1 => lbl2_n_137, A2 => lbl2_n_135, A3 => lbl2_n_128, ZN => lbl2_n_140);
  lbl2_g2837 : NR3D0BWP7T port map(A1 => lbl2_n_138, A2 => lbl2_n_136, A3 => lbl2_n_129, ZN => lbl2_n_139);
  lbl2_g2838 : OAI221D0BWP7T port map(A1 => lbl2_n_122, A2 => position_1(8), B1 => position_1(4), B2 => lbl2_n_123, C => lbl2_n_134, ZN => lbl2_n_138);
  lbl2_g2839 : OAI221D0BWP7T port map(A1 => lbl2_n_122, A2 => position_0(8), B1 => position_0(4), B2 => lbl2_n_123, C => lbl2_n_133, ZN => lbl2_n_137);
  lbl2_g2840 : AO211D0BWP7T port map(A1 => lbl2_n_122, A2 => position_1(8), B => lbl2_n_132, C => lbl2_n_115, Z => lbl2_n_136);
  lbl2_g2841 : AO211D0BWP7T port map(A1 => lbl2_n_122, A2 => position_0(8), B => lbl2_n_131, C => lbl2_n_116, Z => lbl2_n_135);
  lbl2_g2842 : AOI22D0BWP7T port map(A1 => lbl2_n_123, A2 => position_1(4), B1 => lbl2_n_126, B2 => position_1(3), ZN => lbl2_n_134);
  lbl2_g2843 : AOI22D0BWP7T port map(A1 => lbl2_n_123, A2 => position_0(4), B1 => lbl2_n_126, B2 => position_0(3), ZN => lbl2_n_133);
  lbl2_g2844 : NR2D0BWP7T port map(A1 => lbl2_n_126, A2 => position_1(3), ZN => lbl2_n_132);
  lbl2_g2845 : NR2XD0BWP7T port map(A1 => lbl2_n_126, A2 => position_0(3), ZN => lbl2_n_131);
  lbl2_g2846 : XNR2D1BWP7T port map(A1 => lbl2_y_vec(2), A2 => position_1(7), ZN => lbl2_n_130);
  lbl2_g2847 : CKXOR2D1BWP7T port map(A1 => lbl2_y_vec(4), A2 => position_1(9), Z => lbl2_n_129);
  lbl2_g2848 : CKXOR2D1BWP7T port map(A1 => lbl2_y_vec(4), A2 => position_0(9), Z => lbl2_n_128);
  lbl2_g2849 : XNR2D1BWP7T port map(A1 => lbl2_y_vec(2), A2 => position_0(7), ZN => lbl2_n_127);
  lbl2_g2850 : INVD1BWP7T port map(I => lbl2_central_x_vec(7), ZN => lbl2_n_126);
  lbl2_g2851 : MOAI22D1BWP7T port map(A1 => lbl2_n_75, A2 => lbl2_h_count(7), B1 => lbl2_n_75, B2 => lbl2_h_count(7), ZN => lbl2_central_x_vec(7));
  lbl2_g2852 : MAOI22D0BWP7T port map(A1 => lbl2_central_x_vec(6), A2 => position_1(2), B1 => lbl2_central_x_vec(6), B2 => position_1(2), ZN => lbl2_n_125);
  lbl2_g2853 : MAOI22D0BWP7T port map(A1 => lbl2_central_x_vec(6), A2 => position_0(2), B1 => lbl2_central_x_vec(6), B2 => position_0(2), ZN => lbl2_n_124);
  lbl2_g2854 : AO22D0BWP7T port map(A1 => lbl2_n_53, A2 => lbl2_h_count(1), B1 => lbl2_h_count(2), B2 => lbl2_n_156, Z => lbl2_dx(2));
  lbl2_g2855 : AO22D0BWP7T port map(A1 => lbl2_n_53, A2 => lbl2_h_count(2), B1 => lbl2_h_count(3), B2 => lbl2_n_156, Z => lbl2_dx(3));
  lbl2_g2856 : AO22D0BWP7T port map(A1 => lbl2_n_53, A2 => lbl2_v_count(2), B1 => lbl2_v_count(3), B2 => lbl2_n_156, Z => lbl2_dy_vec(3));
  lbl2_g2857 : AO22D0BWP7T port map(A1 => lbl2_n_53, A2 => lbl2_h_count(0), B1 => lbl2_h_count(1), B2 => lbl2_n_156, Z => lbl2_dx(1));
  lbl2_g2858 : AO22D0BWP7T port map(A1 => lbl2_n_53, A2 => lbl2_v_count(1), B1 => lbl2_v_count(2), B2 => lbl2_n_156, Z => lbl2_dy_vec(2));
  lbl2_g2859 : INVD1BWP7T port map(I => lbl2_n_123, ZN => lbl2_central_x_vec(8));
  lbl2_g2861 : AO22D0BWP7T port map(A1 => lbl2_n_53, A2 => lbl2_v_count(0), B1 => lbl2_v_count(1), B2 => lbl2_n_156, Z => lbl2_dy_vec(1));
  lbl2_g2862 : XNR2D1BWP7T port map(A1 => lbl2_n_146, A2 => lbl2_h_count(8), ZN => lbl2_n_123);
  lbl2_g2863 : MOAI22D0BWP7T port map(A1 => lbl2_n_156, A2 => lbl2_v_count(3), B1 => lbl2_n_156, B2 => lbl2_v_count(6), ZN => lbl2_y_vec(2));
  lbl2_g2864 : MOAI22D0BWP7T port map(A1 => lbl2_n_156, A2 => lbl2_v_count(7), B1 => lbl2_n_156, B2 => lbl2_v_count(8), ZN => lbl2_y_vec(4));
  lbl2_g2865 : MAOI22D0BWP7T port map(A1 => lbl2_n_156, A2 => lbl2_v_count(7), B1 => lbl2_n_156, B2 => lbl2_v_count(6), ZN => lbl2_n_122);
  lbl2_g2866 : CKAN2D1BWP7T port map(A1 => lbl2_n_156, A2 => lbl2_v_count(0), Z => lbl2_dy_vec(0));
  lbl2_g2867 : INR2D1BWP7T port map(A1 => lbl2_h_count(0), B1 => lbl2_n_53, ZN => lbl2_dx(0));
  lbl2_g2868 : INVD1BWP7T port map(I => lbl2_n_53, ZN => lbl2_n_156);
  lbl2_g2869 : XNR2D1BWP7T port map(A1 => lbl2_v_count(5), A2 => position_0(6), ZN => lbl2_n_120);
  lbl2_g2870 : XNR2D1BWP7T port map(A1 => lbl2_v_count(4), A2 => position_1(5), ZN => lbl2_n_119);
  lbl2_g2871 : XNR2D1BWP7T port map(A1 => lbl2_v_count(5), A2 => position_1(6), ZN => lbl2_n_118);
  lbl2_g2872 : ND2D1BWP7T port map(A1 => lbl2_n_147, A2 => lbl2_h_count(5), ZN => lbl2_n_146);
  lbl2_g2873 : NR2XD0BWP7T port map(A1 => lbl2_n_158, A2 => game_state(2), ZN => lbl2_n_53);
  lbl2_g2874 : XNR2D1BWP7T port map(A1 => lbl2_v_count(4), A2 => position_0(5), ZN => lbl2_n_117);
  lbl2_g2875 : CKXOR2D1BWP7T port map(A1 => lbl2_h_count(4), A2 => position_0(0), Z => lbl2_n_116);
  lbl2_g2876 : CKXOR2D0BWP7T port map(A1 => lbl2_h_count(4), A2 => position_1(0), Z => lbl2_n_115);
  lbl2_g2877 : MAOI22D0BWP7T port map(A1 => lbl2_central_x_vec(5), A2 => position_1(1), B1 => lbl2_central_x_vec(5), B2 => position_1(1), ZN => lbl2_n_114);
  lbl2_g2878 : MAOI22D0BWP7T port map(A1 => lbl2_central_x_vec(5), A2 => position_0(1), B1 => lbl2_central_x_vec(5), B2 => position_0(1), ZN => lbl2_n_113);
  lbl2_g2879 : MOAI22D1BWP7T port map(A1 => lbl2_central_x_vec(5), A2 => lbl2_h_count(6), B1 => lbl2_central_x_vec(5), B2 => lbl2_h_count(6), ZN => lbl2_central_x_vec(6));
  lbl2_g2880 : AN2D1BWP7T port map(A1 => lbl2_h_count(6), A2 => lbl2_h_count(7), Z => lbl2_n_147);
  lbl2_g2881 : OR2D1BWP7T port map(A1 => game_state(0), A2 => game_state(1), Z => lbl2_n_158);
  lbl2_g2882 : ND2D1BWP7T port map(A1 => lbl2_h_count(5), A2 => lbl2_h_count(6), ZN => lbl2_n_75);
  lbl2_color_reg_0 : DFD0BWP7T port map(CP => CTS_20, D => lbl2_n_103, Q => UNCONNECTED, QN => lbl2_n_108);
  lbl2_color_reg_1 : DFD0BWP7T port map(CP => CTS_20, D => lbl2_n_106, Q => UNCONNECTED0, QN => lbl2_n_110);
  lbl2_color_reg_2 : DFD0BWP7T port map(CP => CTS_20, D => lbl2_n_105, Q => UNCONNECTED1, QN => lbl2_n_111);
  lbl2_color_reg_3 : DFD0BWP7T port map(CP => CTS_20, D => lbl2_n_104, Q => UNCONNECTED2, QN => lbl2_n_109);
  lbl2_h_sync_reg : DFKSND1BWP7T port map(CP => CTS_20, D => lbl2_n_83, Q => UNCONNECTED3, QN => lbl2_n_91, SN => FE_DBTN24_rst);
  lbl2_v_sync_reg : DFKSND0BWP7T port map(CP => CTS_20, D => FE_OFN1_rst, Q => UNCONNECTED4, QN => lbl2_n_100, SN => lbl2_n_92);
  lbl2_g3647 : IINR4D0BWP7T port map(A1 => lbl2_dx(2), A2 => lbl2_dx(3), B1 => lbl2_n_107, B2 => lbl2_n_88, ZN => x_increment);
  lbl2_g3649 : INVD5BWP7T port map(I => lbl2_n_111, ZN => color_out(2));
  lbl2_g3651 : INVD5BWP7T port map(I => lbl2_n_110, ZN => color_out(1));
  lbl2_g3653 : INVD5BWP7T port map(I => lbl2_n_109, ZN => color_out(3));
  lbl2_g3655 : INVD5BWP7T port map(I => lbl2_n_108, ZN => color_out(0));
  lbl2_g3656 : OAI211D1BWP7T port map(A1 => lbl2_n_53, A2 => lbl2_dx(0), B => lbl2_n_102, C => lbl2_dx(1), ZN => lbl2_n_107);
  lbl2_g3657 : AO222D0BWP7T port map(A1 => lbl2_homescreen_color(1), A2 => lbl2_n_98, B1 => lbl2_pixelator_color(1), B2 => lbl2_n_101, C1 => lbl2_sidebar_color(1), C2 => lbl2_n_96, Z => lbl2_n_106);
  lbl2_g3658 : AO222D0BWP7T port map(A1 => lbl2_homescreen_color(2), A2 => lbl2_n_98, B1 => lbl2_pixelator_color(2), B2 => lbl2_n_101, C1 => lbl2_sidebar_color(2), C2 => lbl2_n_96, Z => lbl2_n_105);
  lbl2_g3659 : AO222D0BWP7T port map(A1 => lbl2_homescreen_color(3), A2 => lbl2_n_98, B1 => lbl2_pixelator_color(3), B2 => lbl2_n_101, C1 => lbl2_sidebar_color(3), C2 => lbl2_n_96, Z => lbl2_n_104);
  lbl2_g3660 : AO222D0BWP7T port map(A1 => lbl2_homescreen_color(0), A2 => lbl2_n_98, B1 => lbl2_pixelator_color(0), B2 => lbl2_n_101, C1 => lbl2_sidebar_color(0), C2 => lbl2_n_96, Z => lbl2_n_103);
  lbl2_g3661 : MOAI22D0BWP7T port map(A1 => lbl2_n_99, A2 => lbl2_n_94, B1 => lbl2_n_99, B2 => lbl2_n_94, ZN => lbl2_n_102);
  lbl2_g3662 : INR3D0BWP7T port map(A1 => lbl2_n_69, B1 => lbl2_n_95, B2 => lbl2_n_85, ZN => y_increment);
  lbl2_g3664 : INVD5BWP7T port map(I => lbl2_n_100, ZN => v_sync_out);
  lbl2_g3665 : NR2D1BWP7T port map(A1 => lbl2_n_97, A2 => lbl2_n_53, ZN => lbl2_n_101);
  lbl2_g3666 : INR2XD0BWP7T port map(A1 => lbl2_n_85, B1 => lbl2_n_95, ZN => reset_vga_mem);
  lbl2_g3667 : AOI222D0BWP7T port map(A1 => lbl2_n_53, A2 => lbl2_n_87, B1 => lbl2_n_89, B2 => lbl2_n_73, C1 => lbl2_n_156, C2 => lbl2_h_count(8), ZN => lbl2_n_99);
  lbl2_g3668 : NR2D1BWP7T port map(A1 => lbl2_n_97, A2 => lbl2_n_156, ZN => lbl2_n_98);
  lbl2_g3669 : CKND2D1BWP7T port map(A1 => lbl2_n_93, A2 => lbl2_n_90, ZN => lbl2_n_97);
  lbl2_g3670 : INR2D1BWP7T port map(A1 => lbl2_n_93, B1 => lbl2_n_90, ZN => lbl2_n_96);
  lbl2_g3671 : OR4D1BWP7T port map(A1 => lbl2_h_count(3), A2 => lbl2_n_73, A3 => lbl2_n_78, A4 => lbl2_n_88, Z => lbl2_n_95);
  lbl2_g3672 : AO32D1BWP7T port map(A1 => lbl2_n_53, A2 => lbl2_n_86, A3 => lbl2_n_73, B1 => lbl2_n_156, B2 => lbl2_h_count(9), Z => lbl2_n_94);
  lbl2_g3673 : NR4D0BWP7T port map(A1 => lbl2_n_88, A2 => lbl2_n_79, A3 => lbl2_n_82, A4 => FE_OFN1_rst, ZN => lbl2_n_93);
  lbl2_g3674 : OAI31D0BWP7T port map(A1 => FE_PHN238_lbl2_v_count_9, A2 => lbl2_v_count(4), A3 => lbl2_n_81, B => FE_DBTN24_rst, ZN => lbl2_n_92);
  lbl2_g3676 : INVD5BWP7T port map(I => lbl2_n_91, ZN => h_sync_out);
  lbl2_g3677 : INR3D0BWP7T port map(A1 => lbl2_h_count(6), B1 => lbl2_n_229, B2 => lbl2_n_227, ZN => lbl2_n_89);
  lbl2_g3678 : AOI211XD0BWP7T port map(A1 => lbl2_n_146, A2 => lbl2_n_66, B => lbl2_n_84, C => lbl2_n_68, ZN => lbl2_n_90);
  lbl2_g3679 : OAI21D0BWP7T port map(A1 => lbl2_n_158, A2 => lbl2_n_59, B => busy, ZN => lbl2_n_88);
  lbl2_g3680 : MOAI22D0BWP7T port map(A1 => lbl2_n_75, A2 => lbl2_n_74, B1 => lbl2_n_75, B2 => lbl2_h_count(7), ZN => lbl2_n_87);
  lbl2_g3681 : MOAI22D0BWP7T port map(A1 => lbl2_n_228, A2 => lbl2_h_count(8), B1 => lbl2_n_228, B2 => lbl2_h_count(8), ZN => lbl2_n_86);
  lbl2_g3682 : OAI22D0BWP7T port map(A1 => lbl2_n_70, A2 => lbl2_h_count(5), B1 => lbl2_n_146, B2 => lbl2_n_50, ZN => lbl2_n_84);
  lbl2_g3683 : INR2XD0BWP7T port map(A1 => lbl2_n_77, B1 => FE_PHN238_lbl2_v_count_9, ZN => busy);
  lbl2_g3684 : NR4D0BWP7T port map(A1 => lbl2_n_230, A2 => lbl2_y_vec(4), A3 => lbl2_v_count(4), A4 => lbl2_v_count(5), ZN => lbl2_n_85);
  lbl2_g3685 : AOI21D0BWP7T port map(A1 => lbl2_n_72, A2 => lbl2_n_75, B => FE_OFN1_rst, ZN => lbl2_n_83);
  lbl2_g3686 : OA21D0BWP7T port map(A1 => lbl2_n_71, A2 => lbl2_n_74, B => lbl2_n_68, Z => lbl2_n_82);
  lbl2_g3687 : IIND4D0BWP7T port map(A1 => lbl2_n_77, A2 => lbl2_v_count(2), B1 => lbl2_v_count(3), B2 => lbl2_v_count(1), ZN => lbl2_n_81);
  lbl2_g3689 : AOI211XD0BWP7T port map(A1 => lbl2_n_60, A2 => lbl2_h_count(7), B => lbl2_n_147, C => lbl2_n_67, ZN => lbl2_n_79);
  lbl2_g3690 : OR4D1BWP7T port map(A1 => lbl2_h_count(1), A2 => lbl2_h_count(2), A3 => lbl2_h_count(0), A4 => lbl2_n_71, Z => lbl2_n_78);
  lbl2_g3691 : ND4D0BWP7T port map(A1 => lbl2_v_count(5), A2 => lbl2_v_count(7), A3 => lbl2_v_count(8), A4 => lbl2_v_count(6), ZN => lbl2_n_77);
  lbl2_g3694 : INVD1BWP7T port map(I => lbl2_n_72, ZN => lbl2_n_73);
  lbl2_g3695 : IND2D1BWP7T port map(A1 => lbl2_h_count(7), B1 => lbl2_n_67, ZN => lbl2_n_74);
  lbl2_g3696 : NR2XD0BWP7T port map(A1 => lbl2_n_67, A2 => lbl2_h_count(7), ZN => lbl2_n_72);
  lbl2_g3697 : ND3D0BWP7T port map(A1 => lbl2_central_x_vec(8), A2 => lbl2_central_x_vec(7), A3 => lbl2_central_x_vec(6), ZN => lbl2_n_70);
  lbl2_g3698 : NR4D0BWP7T port map(A1 => lbl2_dy_vec(1), A2 => lbl2_dy_vec(2), A3 => lbl2_dy_vec(3), A4 => lbl2_dy_vec(0), ZN => lbl2_n_69);
  lbl2_g3699 : IND2D1BWP7T port map(A1 => lbl2_h_count(6), B1 => lbl2_n_229, ZN => lbl2_n_71);
  lbl2_g3700 : INVD1BWP7T port map(I => lbl2_n_66, ZN => lbl2_n_67);
  lbl2_g3701 : ND2D0BWP7T port map(A1 => lbl2_h_count(5), A2 => lbl2_h_count(3), ZN => lbl2_n_65);
  lbl2_g3702 : INR2D1BWP7T port map(A1 => lbl2_h_count(8), B1 => lbl2_n_50, ZN => lbl2_n_68);
  lbl2_g3703 : NR2XD0BWP7T port map(A1 => lbl2_h_count(9), A2 => lbl2_h_count(8), ZN => lbl2_n_66);
  lbl2_g3708 : INVD0BWP7T port map(I => lbl2_n_229, ZN => lbl2_n_60);
  lbl2_g3709 : CKND1BWP7T port map(I => game_state(2), ZN => lbl2_n_59);
  lbl2_g2160 : MOAI22D0BWP7T port map(A1 => lbl2_n_51, A2 => lbl2_h_count(5), B1 => lbl2_n_51, B2 => lbl2_h_count(5), ZN => lbl2_n_149);
  lbl2_g2161 : MOAI22D0BWP7T port map(A1 => lbl2_n_52, A2 => lbl2_h_count(6), B1 => lbl2_n_52, B2 => lbl2_h_count(6), ZN => lbl2_n_150);
  lbl2_g2162 : IOA21D1BWP7T port map(A1 => lbl2_h_count(4), A2 => lbl2_h_count(9), B => lbl2_n_51, ZN => lbl2_n_148);
  lbl2_g2163 : AO22D0BWP7T port map(A1 => lbl2_n_50, A2 => direction_between(1), B1 => direction_between(3), B2 => lbl2_h_count(9), Z => lbl2_n_153);
  lbl2_g2164 : NR2D0BWP7T port map(A1 => lbl2_n_229, A2 => lbl2_h_count(9), ZN => lbl2_n_52);
  lbl2_g2165 : AO22D0BWP7T port map(A1 => lbl2_n_50, A2 => direction_between(0), B1 => direction_between(2), B2 => lbl2_h_count(9), Z => lbl2_n_152);
  lbl2_g2166 : AO22D0BWP7T port map(A1 => lbl2_n_50, A2 => boost_audio_0, B1 => boost_audio_1, B2 => lbl2_h_count(9), Z => lbl2_n_154);
  lbl2_g2167 : AO22D0BWP7T port map(A1 => lbl2_n_50, A2 => player_state_0(0), B1 => player_state_1(0), B2 => lbl2_h_count(9), Z => lbl2_n_151);
  lbl2_g2169 : IND2D1BWP7T port map(A1 => lbl2_h_count(4), B1 => lbl2_n_50, ZN => lbl2_n_51);
  lbl2_borders_synced_reg_0 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN68_lbl2_borders_synced_0, DB => borders(0), Q => lbl2_borders_synced(0), SA => FE_OFN0_lbl2_n_2);
  lbl2_borders_synced_reg_1 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN94_lbl2_borders_synced_1, DB => borders(1), Q => lbl2_borders_synced(1), SA => FE_OFN0_lbl2_n_2);
  lbl2_borders_synced_reg_2 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN83_lbl2_borders_synced_2, DB => borders(2), Q => lbl2_borders_synced(2), SA => FE_OFN0_lbl2_n_2);
  lbl2_borders_synced_reg_3 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN73_lbl2_borders_synced_3, DB => borders(3), Q => lbl2_borders_synced(3), SA => FE_OFN0_lbl2_n_2);
  lbl2_borders_synced_reg_4 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN74_lbl2_borders_synced_4, DB => borders(4), Q => lbl2_borders_synced(4), SA => FE_OFN0_lbl2_n_2);
  lbl2_borders_synced_reg_5 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN93_lbl2_borders_synced_5, DB => borders(5), Q => lbl2_borders_synced(5), SA => FE_OFN0_lbl2_n_2);
  lbl2_borders_synced_reg_6 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN85_lbl2_borders_synced_6, DB => borders(6), Q => lbl2_borders_synced(6), SA => FE_OFN0_lbl2_n_2);
  lbl2_borders_synced_reg_7 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN82_lbl2_borders_synced_7, DB => borders(7), Q => lbl2_borders_synced(7), SA => FE_OFN0_lbl2_n_2);
  lbl2_data_synced_reg_0 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN116_lbl2_data_synced_0, DB => FE_PHN217_read_memory_in_0, Q => lbl2_data_synced(0), SA => FE_OFN0_lbl2_n_2);
  lbl2_data_synced_reg_1 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN129_lbl2_data_synced_1, DB => FE_PHN205_read_memory_in_1, Q => lbl2_data_synced(1), SA => FE_OFN0_lbl2_n_2);
  lbl2_data_synced_reg_2 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN133_lbl2_data_synced_2, DB => FE_PHN201_read_memory_in_2, Q => lbl2_data_synced(2), SA => FE_OFN0_lbl2_n_2);
  lbl2_data_synced_reg_3 : DFXQD1BWP7T port map(CP => CTS_20, DA => FE_PHN101_lbl2_data_synced_3, DB => FE_PHN153_read_memory_in_3, Q => lbl2_data_synced(3), SA => FE_OFN0_lbl2_n_2);
  lbl2_data_synced_reg_4 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN109_lbl2_data_synced_4, DB => FE_PHN235_read_memory_in_4, Q => lbl2_data_synced(4), SA => FE_OFN0_lbl2_n_2);
  lbl2_data_synced_reg_5 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN122_lbl2_data_synced_5, DB => FE_PHN231_read_memory_in_5, Q => lbl2_data_synced(5), SA => FE_OFN0_lbl2_n_2);
  lbl2_data_synced_reg_6 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN120_lbl2_data_synced_6, DB => FE_PHN198_read_memory_in_6, Q => lbl2_data_synced(6), SA => FE_OFN0_lbl2_n_2);
  lbl2_data_synced_reg_7 : DFXQD1BWP7T port map(CP => CTS_20, DA => FE_PHN79_lbl2_data_synced_7, DB => FE_PHN193_read_memory_in_7, Q => lbl2_data_synced(7), SA => FE_OFN0_lbl2_n_2);
  lbl2_h_count_reg_0 : DFKCNQD1BWP7T port map(CN => FE_PHN229_lbl2_n_21, CP => CTS_20, D => lbl2_n_9, Q => lbl2_h_count(0));
  lbl2_h_count_reg_1 : DFKCNQD1BWP7T port map(CN => lbl2_n_9, CP => CTS_20, D => lbl2_n_25, Q => lbl2_h_count(1));
  lbl2_h_count_reg_2 : DFKCNQD1BWP7T port map(CN => lbl2_n_9, CP => CTS_20, D => lbl2_n_28, Q => lbl2_h_count(2));
  lbl2_h_count_reg_3 : DFKCNQD1BWP7T port map(CN => lbl2_n_9, CP => CTS_20, D => lbl2_n_31, Q => lbl2_h_count(3));
  lbl2_h_count_reg_4 : DFKCNQD1BWP7T port map(CN => lbl2_n_9, CP => CTS_20, D => lbl2_n_34, Q => lbl2_h_count(4));
  lbl2_h_count_reg_6 : DFKCNQD1BWP7T port map(CN => lbl2_n_9, CP => CTS_21, D => lbl2_n_40, Q => lbl2_h_count(6));
  lbl2_h_count_reg_7 : DFKCNQD1BWP7T port map(CN => lbl2_n_9, CP => CTS_20, D => lbl2_n_43, Q => lbl2_h_count(7));
  lbl2_h_count_reg_8 : DFKCNQD1BWP7T port map(CN => lbl2_n_9, CP => CTS_20, D => lbl2_n_46, Q => lbl2_h_count(8));
  lbl2_jumps_synced_reg_0 : DFXQD1BWP7T port map(CP => CTS_21, DA => FE_PHN75_lbl2_jumps_synced_0, DB => ramps(0), Q => lbl2_jumps_synced(0), SA => FE_OFN0_lbl2_n_2);
  lbl2_jumps_synced_reg_1 : DFXQD1BWP7T port map(CP => CTS_21, DA => FE_PHN71_lbl2_jumps_synced_1, DB => ramps(1), Q => lbl2_jumps_synced(1), SA => FE_OFN0_lbl2_n_2);
  lbl2_jumps_synced_reg_2 : DFXQD1BWP7T port map(CP => CTS_21, DA => FE_PHN67_lbl2_jumps_synced_2, DB => ramps(2), Q => lbl2_jumps_synced(2), SA => FE_OFN0_lbl2_n_2);
  lbl2_jumps_synced_reg_3 : DFXQD1BWP7T port map(CP => CTS_18, DA => FE_PHN77_lbl2_jumps_synced_3, DB => ramps(3), Q => lbl2_jumps_synced(3), SA => FE_OFN0_lbl2_n_2);
  lbl2_jumps_synced_reg_4 : DFXQD1BWP7T port map(CP => CTS_21, DA => FE_PHN69_lbl2_jumps_synced_4, DB => ramps(4), Q => lbl2_jumps_synced(4), SA => FE_OFN0_lbl2_n_2);
  lbl2_jumps_synced_reg_5 : DFXQD1BWP7T port map(CP => CTS_21, DA => FE_PHN78_lbl2_jumps_synced_5, DB => ramps(5), Q => lbl2_jumps_synced(5), SA => FE_OFN0_lbl2_n_2);
  lbl2_jumps_synced_reg_6 : DFXQD1BWP7T port map(CP => CTS_21, DA => FE_PHN76_lbl2_jumps_synced_6, DB => ramps(6), Q => lbl2_jumps_synced(6), SA => FE_OFN0_lbl2_n_2);
  lbl2_jumps_synced_reg_7 : DFXQD1BWP7T port map(CP => CTS_21, DA => FE_PHN323_lbl2_jumps_synced_7, DB => ramps(7), Q => lbl2_jumps_synced(7), SA => FE_OFN0_lbl2_n_2);
  lbl2_v_count_reg_0 : DFQD1BWP7T port map(CP => CTS_20, D => lbl2_n_23, Q => lbl2_v_count(0));
  lbl2_v_count_reg_1 : DFQD1BWP7T port map(CP => CTS_20, D => lbl2_n_26, Q => lbl2_v_count(1));
  lbl2_v_count_reg_2 : DFQD1BWP7T port map(CP => CTS_20, D => lbl2_n_29, Q => lbl2_v_count(2));
  lbl2_v_count_reg_3 : DFQD1BWP7T port map(CP => CTS_20, D => lbl2_n_32, Q => lbl2_v_count(3));
  lbl2_v_count_reg_4 : DFQD1BWP7T port map(CP => CTS_20, D => lbl2_n_35, Q => lbl2_v_count(4));
  lbl2_v_count_reg_5 : DFQD1BWP7T port map(CP => CTS_21, D => lbl2_n_38, Q => lbl2_v_count(5));
  lbl2_v_count_reg_6 : DFQD1BWP7T port map(CP => CTS_21, D => lbl2_n_41, Q => lbl2_v_count(6));
  lbl2_v_count_reg_7 : DFQD1BWP7T port map(CP => CTS_20, D => lbl2_n_44, Q => lbl2_v_count(7));
  lbl2_v_count_reg_8 : DFQD1BWP7T port map(CP => CTS_20, D => lbl2_n_47, Q => lbl2_v_count(8));
  lbl2_v_count_reg_9 : DFQD1BWP7T port map(CP => CTS_20, D => lbl2_n_49, Q => lbl2_v_count(9));
  lbl2_g3249 : AO22D0BWP7T port map(A1 => lbl2_n_48, A2 => lbl2_n_20, B1 => FE_PHN316_lbl2_v_count_9, B2 => lbl2_n_9, Z => lbl2_n_49);
  lbl2_g3252 : AO22D0BWP7T port map(A1 => lbl2_n_46, A2 => lbl2_n_20, B1 => FE_PHN150_lbl2_v_count_8, B2 => lbl2_n_9, Z => lbl2_n_47);
  lbl2_g3253 : MOAI22D0BWP7T port map(A1 => lbl2_n_45, A2 => lbl2_n_15, B1 => lbl2_n_45, B2 => lbl2_n_15, ZN => lbl2_n_48);
  lbl2_g3254 : HA1D0BWP7T port map(A => lbl2_n_11, B => lbl2_n_42, CO => lbl2_n_45, S => lbl2_n_46);
  lbl2_g3257 : AO22D0BWP7T port map(A1 => lbl2_n_43, A2 => lbl2_n_20, B1 => FE_PHN336_lbl2_v_count_7, B2 => lbl2_n_9, Z => lbl2_n_44);
  lbl2_g3258 : HA1D0BWP7T port map(A => lbl2_n_16, B => lbl2_n_39, CO => lbl2_n_42, S => lbl2_n_43);
  lbl2_g3261 : AO22D0BWP7T port map(A1 => lbl2_n_40, A2 => lbl2_n_20, B1 => FE_PHN138_lbl2_v_count_6, B2 => lbl2_n_9, Z => lbl2_n_41);
  lbl2_g3262 : HA1D0BWP7T port map(A => lbl2_n_18, B => lbl2_n_36, CO => lbl2_n_39, S => lbl2_n_40);
  lbl2_g3265 : AO22D0BWP7T port map(A1 => lbl2_n_37, A2 => lbl2_n_20, B1 => lbl2_v_count(5), B2 => lbl2_n_9, Z => lbl2_n_38);
  lbl2_g3266 : HA1D0BWP7T port map(A => lbl2_n_17, B => lbl2_n_33, CO => lbl2_n_36, S => lbl2_n_37);
  lbl2_g3269 : AO22D0BWP7T port map(A1 => lbl2_n_34, A2 => lbl2_n_20, B1 => lbl2_v_count(4), B2 => lbl2_n_9, Z => lbl2_n_35);
  lbl2_g3270 : HA1D0BWP7T port map(A => lbl2_n_12, B => lbl2_n_30, CO => lbl2_n_33, S => lbl2_n_34);
  lbl2_g3273 : AO22D0BWP7T port map(A1 => lbl2_n_31, A2 => lbl2_n_20, B1 => lbl2_v_count(3), B2 => lbl2_n_9, Z => lbl2_n_32);
  lbl2_g3274 : HA1D0BWP7T port map(A => lbl2_n_13, B => lbl2_n_27, CO => lbl2_n_30, S => lbl2_n_31);
  lbl2_g3277 : AO22D0BWP7T port map(A1 => lbl2_n_28, A2 => lbl2_n_20, B1 => lbl2_v_count(2), B2 => lbl2_n_9, Z => lbl2_n_29);
  lbl2_g3278 : HA1D0BWP7T port map(A => lbl2_n_14, B => lbl2_n_24, CO => lbl2_n_27, S => lbl2_n_28);
  lbl2_g3281 : AO22D0BWP7T port map(A1 => lbl2_n_25, A2 => lbl2_n_20, B1 => lbl2_v_count(1), B2 => lbl2_n_9, Z => lbl2_n_26);
  lbl2_g3282 : HA1D0BWP7T port map(A => lbl2_n_22, B => lbl2_n_10, CO => lbl2_n_24, S => lbl2_n_25);
  lbl2_g3285 : MOAI22D0BWP7T port map(A1 => lbl2_n_19, A2 => lbl2_n_22, B1 => lbl2_n_9, B2 => lbl2_v_count(0), ZN => lbl2_n_23);
  lbl2_g3286 : INVD0BWP7T port map(I => lbl2_n_21, ZN => lbl2_n_22);
  lbl2_g3287 : INVD0BWP7T port map(I => lbl2_n_20, ZN => lbl2_n_19);
  lbl2_g3288 : AO21D0BWP7T port map(A1 => lbl2_n_7, A2 => lbl2_v_count(6), B => lbl2_h_count(6), Z => lbl2_n_18);
  lbl2_g3289 : AO21D0BWP7T port map(A1 => lbl2_n_7, A2 => lbl2_v_count(5), B => lbl2_h_count(5), Z => lbl2_n_17);
  lbl2_g3290 : AO21D0BWP7T port map(A1 => lbl2_n_7, A2 => lbl2_v_count(7), B => lbl2_h_count(7), Z => lbl2_n_16);
  lbl2_g3291 : AOI22D0BWP7T port map(A1 => lbl2_n_7, A2 => lbl2_v_count(0), B1 => lbl2_n_8, B2 => lbl2_h_count(0), ZN => lbl2_n_21);
  lbl2_g3292 : AOI211XD0BWP7T port map(A1 => lbl2_n_6, A2 => FE_PHN238_lbl2_v_count_9, B => lbl2_n_8, C => FE_OFN1_rst, ZN => lbl2_n_20);
  lbl2_g3293 : AOI22D0BWP7T port map(A1 => lbl2_n_7, A2 => FE_PHN238_lbl2_v_count_9, B1 => lbl2_n_8, B2 => lbl2_h_count(9), ZN => lbl2_n_15);
  lbl2_g3294 : AO22D0BWP7T port map(A1 => lbl2_n_7, A2 => lbl2_v_count(2), B1 => lbl2_h_count(2), B2 => lbl2_n_8, Z => lbl2_n_14);
  lbl2_g3295 : AO22D0BWP7T port map(A1 => lbl2_n_7, A2 => lbl2_v_count(3), B1 => lbl2_h_count(3), B2 => lbl2_n_8, Z => lbl2_n_13);
  lbl2_g3296 : AO22D0BWP7T port map(A1 => lbl2_n_7, A2 => lbl2_v_count(4), B1 => lbl2_h_count(4), B2 => lbl2_n_8, Z => lbl2_n_12);
  lbl2_g3297 : AO22D0BWP7T port map(A1 => lbl2_n_7, A2 => lbl2_v_count(8), B1 => lbl2_h_count(8), B2 => lbl2_n_8, Z => lbl2_n_11);
  lbl2_g3298 : AO22D0BWP7T port map(A1 => lbl2_n_7, A2 => lbl2_v_count(1), B1 => lbl2_h_count(1), B2 => lbl2_n_8, Z => lbl2_n_10);
  lbl2_g3299 : NR2XD0BWP7T port map(A1 => lbl2_n_7, A2 => FE_OFN1_rst, ZN => lbl2_n_9);
  lbl2_g3300 : INVD1BWP7T port map(I => lbl2_n_8, ZN => lbl2_n_7);
  lbl2_g3301 : IND4D0BWP7T port map(A1 => lbl2_h_count(7), B1 => lbl2_h_count(8), B2 => lbl2_h_count(9), B3 => lbl2_n_5, ZN => lbl2_n_8);
  lbl2_g3302 : INR4D0BWP7T port map(A1 => lbl2_n_4, B1 => lbl2_v_count(8), B2 => lbl2_v_count(7), B3 => lbl2_v_count(6), ZN => lbl2_n_6);
  lbl2_g3315 : INR4D0BWP7T port map(A1 => lbl2_h_count(4), B1 => lbl2_h_count(6), B2 => lbl2_h_count(5), B3 => lbl2_n_1, ZN => lbl2_n_5);
  lbl2_g3328 : NR3D0BWP7T port map(A1 => lbl2_n_3, A2 => lbl2_v_count(5), A3 => lbl2_v_count(4), ZN => lbl2_n_4);
  lbl2_g3329 : IIND4D0BWP7T port map(A1 => lbl2_v_count(0), A2 => lbl2_v_count(1), B1 => lbl2_v_count(2), B2 => lbl2_v_count(3), ZN => lbl2_n_3);
  lbl2_g3330 : ND4D0BWP7T port map(A1 => lbl2_h_count(0), A2 => lbl2_h_count(2), A3 => lbl2_h_count(1), A4 => lbl2_h_count(3), ZN => lbl2_n_1);
  lbl2_g3331 : ND4D0BWP7T port map(A1 => lbl2_n_0, A2 => lbl2_dx(1), A3 => lbl2_dx(3), A4 => lbl2_dx(2), ZN => lbl2_n_2);
  lbl2_g3332 : IND2D1BWP7T port map(A1 => lbl2_dx(0), B1 => lbl2_n_156, ZN => lbl2_n_0);
  lbl2_g2 : AOI22D0BWP7T port map(A1 => lbl2_n_53, A2 => lbl2_n_65, B1 => lbl2_n_156, B2 => lbl2_h_count(7), ZN => lbl2_n_227);
  lbl2_g3717 : INR2D1BWP7T port map(A1 => lbl2_h_count(3), B1 => lbl2_n_146, ZN => lbl2_n_228);
  lbl2_g3718 : NR2XD0BWP7T port map(A1 => lbl2_h_count(5), A2 => lbl2_h_count(4), ZN => lbl2_n_229);
  lbl2_h_count_reg_5 : DFKCND1BWP7T port map(CN => lbl2_n_9, CP => CTS_21, D => lbl2_n_37, Q => lbl2_h_count(5), QN => lbl2_central_x_vec(5));
  lbl2_h_count_reg_9 : DFKCND1BWP7T port map(CN => lbl2_n_9, CP => CTS_20, D => lbl2_n_48, Q => lbl2_h_count(9), QN => lbl2_n_50);
  lbl2_g3723 : IND2D1BWP7T port map(A1 => lbl2_y_vec(2), B1 => lbl2_n_122, ZN => lbl2_n_230);
  lbl3_dir_out_reg_3 : DFKCNQD1BWP7T port map(CN => lbl3_temp1(3), CP => CTS_20, D => FE_DBTN24_rst, Q => direction_between(3));
  lbl3_dir_out_reg_2 : DFKCNQD1BWP7T port map(CN => lbl3_temp1(2), CP => CTS_20, D => FE_DBTN24_rst, Q => direction_between(2));
  lbl3_dir_out_reg_0 : DFKCNQD1BWP7T port map(CN => FE_PHN48_lbl3_temp1_0, CP => CTS_20, D => FE_DBTN24_rst, Q => direction_between(0));
  lbl3_start_out_reg : DFKCNQD1BWP7T port map(CN => FE_PHN50_lbl3_temp2, CP => CTS_20, D => FE_DBTN24_rst, Q => start_between);
  lbl3_dir_out_reg_1 : DFKCNQD1BWP7T port map(CN => FE_PHN55_lbl3_temp1_1, CP => CTS_20, D => FE_DBTN24_rst, Q => direction_between(1));
  lbl3_temp1_reg_1 : DFKCNQD1BWP7T port map(CN => FE_PHN127_direction_in_1, CP => CTS_20, D => FE_DBTN24_rst, Q => lbl3_temp1(1));
  lbl3_temp1_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN328_direction_in_2, CP => CTS_20, D => FE_DBTN24_rst, Q => FE_PHN29_lbl3_temp1_2);
  lbl3_temp1_reg_3 : DFKCNQD1BWP7T port map(CN => FE_PHN103_direction_in_3, CP => CTS_20, D => FE_DBTN24_rst, Q => FE_PHN32_lbl3_temp1_3);
  lbl3_temp2_reg : DFKCNQD1BWP7T port map(CN => FE_PHN65_start_in, CP => CTS_20, D => FE_DBTN24_rst, Q => lbl3_temp2);
  lbl3_temp1_reg_0 : DFKCNQD1BWP7T port map(CN => FE_PHN134_direction_in_0, CP => CTS_20, D => FE_DBTN24_rst, Q => lbl3_temp1(0));
  lbl2_dec0_g100 : AO22D0BWP7T port map(A1 => lbl2_dec0_n_2, A2 => lbl2_data_synced(0), B1 => lbl2_data_synced(1), B2 => lbl2_dec0_n_1, Z => lbl2_walls(2));
  lbl2_dec0_g101 : IOA21D1BWP7T port map(A1 => lbl2_dec0_n_2, A2 => lbl2_dec0_n_0, B => lbl2_dec0_n_5, ZN => lbl2_walls(0));
  lbl2_dec0_g102 : IND2D1BWP7T port map(A1 => lbl2_dec0_n_2, B1 => lbl2_dec0_n_3, ZN => lbl2_walls(1));
  lbl2_dec0_g103 : IOA21D1BWP7T port map(A1 => lbl2_dec0_n_0, A2 => lbl2_data_synced(2), B => lbl2_data_synced(1), ZN => lbl2_dec0_n_5);
  lbl2_dec0_g104 : IOA21D1BWP7T port map(A1 => lbl2_data_synced(1), A2 => lbl2_data_synced(2), B => lbl2_dec0_n_3, ZN => lbl2_walls(3));
  lbl2_dec0_g105 : IND2D1BWP7T port map(A1 => lbl2_data_synced(2), B1 => lbl2_data_synced(0), ZN => lbl2_dec0_n_3);
  lbl2_dec0_g106 : ND2D0BWP7T port map(A1 => lbl2_data_synced(0), A2 => lbl2_data_synced(2), ZN => lbl2_dec0_n_1);
  lbl2_dec0_g107 : INR2D1BWP7T port map(A1 => lbl2_data_synced(2), B1 => lbl2_data_synced(1), ZN => lbl2_dec0_n_2);
  lbl2_dec0_g108 : CKND1BWP7T port map(I => lbl2_data_synced(0), ZN => lbl2_dec0_n_0);
  lbl4_g7892 : IND2D1BWP7T port map(A1 => lbl4_n_86, B1 => lbl4_n_147, ZN => borders(4));
  lbl4_g7893 : IND3D1BWP7T port map(A1 => ramps(5), B1 => lbl4_n_111, B2 => lbl4_n_138, ZN => borders(1));
  lbl4_g7894 : IND2D1BWP7T port map(A1 => ramps(4), B1 => lbl4_n_142, ZN => borders(0));
  lbl4_g7895 : IND4D0BWP7T port map(A1 => lbl4_n_123, B1 => lbl4_n_115, B2 => lbl4_n_126, B3 => lbl4_n_141, ZN => borders(7));
  lbl4_g7896 : AOI221D0BWP7T port map(A1 => lbl4_n_134, A2 => lbl4_n_29, B1 => lbl4_n_97, B2 => lbl4_n_44, C => ramps(0), ZN => lbl4_n_147);
  lbl4_g7897 : IND3D1BWP7T port map(A1 => ramps(7), B1 => lbl4_n_127, B2 => lbl4_n_137, ZN => borders(3));
  lbl4_g7898 : AO221D0BWP7T port map(A1 => lbl4_n_134, A2 => lbl4_n_12, B1 => lbl4_n_95, B2 => lbl4_n_29, C => ramps(2), Z => borders(6));
  lbl4_g7899 : ND3D0BWP7T port map(A1 => lbl4_n_140, A2 => lbl4_n_120, A3 => lbl4_n_124, ZN => borders(5));
  lbl4_g7900 : AO211D0BWP7T port map(A1 => lbl4_n_110, A2 => lbl4_n_41, B => lbl4_n_130, C => ramps(6), Z => borders(2));
  lbl4_g7901 : AOI221D0BWP7T port map(A1 => lbl4_n_122, A2 => lbl4_n_29, B1 => lbl4_n_97, B2 => lbl4_n_80, C => lbl4_n_86, ZN => lbl4_n_142);
  lbl4_g7902 : AOI32D1BWP7T port map(A1 => lbl4_n_114, A2 => lbl4_n_9, A3 => lbl4_n_2, B1 => lbl4_n_104, B2 => lbl4_n_106, ZN => lbl4_n_141);
  lbl4_g7903 : AOI33D1BWP7T port map(A1 => lbl4_n_114, A2 => x_address(0), A3 => lbl4_n_2, B1 => lbl4_n_106, B2 => lbl4_n_76, B3 => start_position_0(3), ZN => lbl4_n_140);
  lbl4_g7904 : AOI33D1BWP7T port map(A1 => lbl4_n_112, A2 => x_address(0), A3 => lbl4_n_2, B1 => lbl4_n_105, B2 => lbl4_n_76, B3 => start_position_0(3), ZN => lbl4_n_138);
  lbl4_g7905 : AOI32D1BWP7T port map(A1 => lbl4_n_112, A2 => lbl4_n_9, A3 => lbl4_n_2, B1 => lbl4_n_104, B2 => lbl4_n_105, ZN => lbl4_n_137);
  lbl4_g7906 : OAI33D1BWP7T port map(A1 => lbl4_n_13, A2 => lbl4_n_37, A3 => lbl4_n_118, B1 => lbl4_n_42, B2 => lbl4_n_48, B3 => lbl4_n_67, ZN => ramps(2));
  lbl4_g7907 : OAI31D1BWP7T port map(A1 => y_address(4), A2 => lbl4_n_19, A3 => lbl4_n_92, B => lbl4_n_119, ZN => ramps(5));
  lbl4_g7908 : OAI31D1BWP7T port map(A1 => lbl4_n_19, A2 => lbl4_n_61, A3 => lbl4_n_84, B => lbl4_n_121, ZN => ramps(7));
  lbl4_g7909 : OAI31D0BWP7T port map(A1 => y_address(2), A2 => lbl4_n_46, A3 => lbl4_n_85, B => lbl4_n_125, ZN => lbl4_n_134);
  lbl4_g7910 : OAI31D1BWP7T port map(A1 => lbl4_n_31, A2 => lbl4_n_54, A3 => lbl4_n_84, B => lbl4_n_124, ZN => ramps(1));
  lbl4_g7911 : AO21D0BWP7T port map(A1 => lbl4_n_98, A2 => lbl4_n_22, B => lbl4_n_123, Z => ramps(3));
  lbl4_g7912 : MOAI22D0BWP7T port map(A1 => lbl4_n_103, A2 => lbl4_n_30, B1 => lbl4_n_117, B2 => lbl4_n_12, ZN => lbl4_n_130);
  lbl4_g7913 : OAI32D1BWP7T port map(A1 => lbl4_n_30, A2 => lbl4_n_67, A3 => lbl4_n_75, B1 => lbl4_n_64, B2 => lbl4_n_118, ZN => ramps(4));
  lbl4_g7914 : AOI31D0BWP7T port map(A1 => lbl4_n_32, A2 => lbl4_n_22, A3 => x_address(2), B => lbl4_n_116, ZN => lbl4_n_127);
  lbl4_g7915 : ND3D0BWP7T port map(A1 => lbl4_n_102, A2 => lbl4_n_22, A3 => x_address(2), ZN => lbl4_n_126);
  lbl4_g7916 : OA31D1BWP7T port map(A1 => lbl4_n_13, A2 => lbl4_n_35, A3 => lbl4_n_90, B => lbl4_n_109, Z => lbl4_n_125);
  lbl4_g7917 : INR2D1BWP7T port map(A1 => lbl4_n_113, B1 => lbl4_n_37, ZN => ramps(6));
  lbl4_g7918 : INR2D1BWP7T port map(A1 => lbl4_n_113, B1 => lbl4_n_38, ZN => ramps(0));
  lbl4_g7919 : AO21D0BWP7T port map(A1 => lbl4_n_110, A2 => lbl4_n_8, B => lbl4_n_117, Z => lbl4_n_122);
  lbl4_g7920 : AOI32D1BWP7T port map(A1 => lbl4_n_89, A2 => lbl4_n_73, A3 => x_address(0), B1 => lbl4_n_93, B2 => lbl4_n_16, ZN => lbl4_n_121);
  lbl4_g7921 : OA32D1BWP7T port map(A1 => lbl4_n_12, A2 => lbl4_n_75, A3 => lbl4_n_77, B1 => lbl4_n_54, B2 => lbl4_n_107, Z => lbl4_n_120);
  lbl4_g7922 : AOI32D1BWP7T port map(A1 => lbl4_n_89, A2 => lbl4_n_53, A3 => lbl4_n_32, B1 => lbl4_n_98, B2 => lbl4_n_16, ZN => lbl4_n_119);
  lbl4_g7923 : OA32D1BWP7T port map(A1 => lbl4_n_15, A2 => lbl4_n_61, A3 => lbl4_n_88, B1 => lbl4_n_19, B2 => lbl4_n_94, Z => lbl4_n_124);
  lbl4_g7924 : OAI33D1BWP7T port map(A1 => lbl4_n_19, A2 => lbl4_n_56, A3 => lbl4_n_88, B1 => y_address(4), B2 => lbl4_n_15, B3 => lbl4_n_92, ZN => lbl4_n_123);
  lbl4_g7925 : NR4D0BWP7T port map(A1 => lbl4_n_79, A2 => lbl4_n_81, A3 => lbl4_n_24, A4 => lbl4_n_9, ZN => lbl4_n_116);
  lbl4_g7926 : OR4XD1BWP7T port map(A1 => lbl4_n_9, A2 => lbl4_n_12, A3 => lbl4_n_75, A4 => lbl4_n_81, Z => lbl4_n_115);
  lbl4_g7927 : AOI21D0BWP7T port map(A1 => lbl4_n_87, A2 => lbl4_n_2, B => lbl4_n_99, ZN => lbl4_n_118);
  lbl4_g7928 : MOAI22D0BWP7T port map(A1 => lbl4_n_96, A2 => lbl4_n_13, B1 => lbl4_n_101, B2 => lbl4_n_44, ZN => lbl4_n_117);
  lbl4_g7929 : AOI21D0BWP7T port map(A1 => lbl4_n_53, A2 => lbl4_n_23, B => lbl4_n_108, ZN => lbl4_n_111);
  lbl4_g7930 : OAI22D0BWP7T port map(A1 => lbl4_n_91, A2 => lbl4_n_43, B1 => lbl4_n_83, B2 => lbl4_n_28, ZN => lbl4_n_114);
  lbl4_g7931 : OAI32D1BWP7T port map(A1 => map_selected(1), A2 => lbl4_n_28, A3 => lbl4_n_82, B1 => lbl4_n_39, B2 => lbl4_n_100, ZN => lbl4_n_113);
  lbl4_g7932 : OAI32D1BWP7T port map(A1 => lbl4_n_28, A2 => lbl4_n_43, A3 => lbl4_n_66, B1 => lbl4_n_72, B2 => lbl4_n_91, ZN => lbl4_n_112);
  lbl4_g7933 : IOA21D1BWP7T port map(A1 => lbl4_n_72, A2 => lbl4_n_43, B => lbl4_n_101, ZN => lbl4_n_109);
  lbl4_g7934 : NR3D0BWP7T port map(A1 => lbl4_n_77, A2 => lbl4_n_79, A3 => lbl4_n_24, ZN => lbl4_n_108);
  lbl4_g7935 : IAO21D0BWP7T port map(A1 => lbl4_n_84, A2 => x_address(4), B => lbl4_n_23, ZN => lbl4_n_107);
  lbl4_g7936 : NR2D0BWP7T port map(A1 => lbl4_n_90, A2 => lbl4_n_58, ZN => lbl4_n_110);
  lbl4_g7937 : AOI21D0BWP7T port map(A1 => lbl4_n_80, A2 => lbl4_n_71, B => lbl4_n_62, ZN => lbl4_n_103);
  lbl4_g7938 : OAI21D0BWP7T port map(A1 => lbl4_n_84, A2 => lbl4_n_7, B => lbl4_n_33, ZN => lbl4_n_102);
  lbl4_g7939 : OAI32D1BWP7T port map(A1 => y_address(3), A2 => lbl4_n_39, A3 => lbl4_n_45, B1 => y_address(4), B2 => lbl4_n_78, ZN => lbl4_n_106);
  lbl4_g7940 : OAI22D0BWP7T port map(A1 => lbl4_n_78, A2 => lbl4_n_5, B1 => lbl4_n_66, B2 => y_address(3), ZN => lbl4_n_105);
  lbl4_g7941 : AOI211D1BWP7T port map(A1 => lbl4_n_70, A2 => lbl4_n_49, B => lbl4_n_10, C => lbl4_n_9, ZN => lbl4_n_104);
  lbl4_g7942 : INVD0BWP7T port map(I => lbl4_n_99, ZN => lbl4_n_100);
  lbl4_g7943 : IND3D0BWP7T port map(A1 => lbl4_n_46, B1 => lbl4_n_34, B2 => lbl4_n_74, ZN => lbl4_n_96);
  lbl4_g7944 : AO21D0BWP7T port map(A1 => lbl4_n_71, A2 => lbl4_n_44, B => lbl4_n_62, Z => lbl4_n_95);
  lbl4_g7945 : OAI21D0BWP7T port map(A1 => lbl4_n_68, A2 => y_address(2), B => lbl4_n_69, ZN => lbl4_n_101);
  lbl4_g7946 : AOI211D0BWP7T port map(A1 => lbl4_n_49, A2 => lbl4_n_57, B => lbl4_n_10, C => FE_PHN247_y_address_3, ZN => lbl4_n_99);
  lbl4_g7947 : NR2D0BWP7T port map(A1 => lbl4_n_84, A2 => lbl4_n_56, ZN => lbl4_n_98);
  lbl4_g7948 : INR3D0BWP7T port map(A1 => lbl4_n_71, B1 => y_address(2), B2 => lbl4_n_37, ZN => lbl4_n_97);
  lbl4_g7949 : INVD0BWP7T port map(I => lbl4_n_93, ZN => lbl4_n_94);
  lbl4_g7950 : INVD0BWP7T port map(I => lbl4_n_89, ZN => lbl4_n_88);
  lbl4_g7951 : NR3D0BWP7T port map(A1 => lbl4_n_65, A2 => lbl4_n_33, A3 => lbl4_n_28, ZN => lbl4_n_87);
  lbl4_g7952 : AOI21D0BWP7T port map(A1 => lbl4_n_47, A2 => lbl4_n_30, B => lbl4_n_85, ZN => lbl4_n_93);
  lbl4_g7953 : OAI211D1BWP7T port map(A1 => lbl4_n_8, A2 => lbl4_n_12, B => lbl4_n_74, C => lbl4_n_34, ZN => lbl4_n_92);
  lbl4_g7954 : OA32D1BWP7T port map(A1 => lbl4_n_5, A2 => lbl4_n_35, A3 => lbl4_n_42, B1 => lbl4_n_28, B2 => lbl4_n_64, Z => lbl4_n_91);
  lbl4_g7955 : AOI32D1BWP7T port map(A1 => lbl4_n_53, A2 => lbl4_n_36, A3 => lbl4_n_2, B1 => lbl4_n_74, B2 => lbl4_n_18, ZN => lbl4_n_90);
  lbl4_g7956 : OAI22D0BWP7T port map(A1 => lbl4_n_68, A2 => lbl4_n_42, B1 => lbl4_n_69, B2 => lbl4_n_12, ZN => lbl4_n_89);
  lbl4_g7957 : IND2D1BWP7T port map(A1 => lbl4_n_66, B1 => lbl4_n_73, ZN => lbl4_n_83);
  lbl4_g7958 : OAI211D1BWP7T port map(A1 => lbl4_n_3, A2 => lbl4_n_20, B => lbl4_n_23, C => lbl4_n_14, ZN => lbl4_n_82);
  lbl4_g7959 : NR3D0BWP7T port map(A1 => lbl4_n_42, A2 => y_address(4), A3 => y_address(3), ZN => lbl4_n_86);
  lbl4_g7960 : IND2D1BWP7T port map(A1 => lbl4_n_58, B1 => lbl4_n_74, ZN => lbl4_n_85);
  lbl4_g7961 : IND2D1BWP7T port map(A1 => lbl4_n_47, B1 => lbl4_n_71, ZN => lbl4_n_84);
  lbl4_g7962 : AOI21D0BWP7T port map(A1 => lbl4_n_59, A2 => x_address(1), B => lbl4_n_50, ZN => lbl4_n_81);
  lbl4_g7963 : OAI21D0BWP7T port map(A1 => lbl4_n_56, A2 => x_address(1), B => lbl4_n_51, ZN => lbl4_n_80);
  lbl4_g7964 : AOI32D1BWP7T port map(A1 => lbl4_n_34, A2 => y_address(2), A3 => y_address(1), B1 => lbl4_n_41, B2 => lbl4_n_27, ZN => lbl4_n_79);
  lbl4_g7965 : AOI22D0BWP7T port map(A1 => lbl4_n_41, A2 => y_address(3), B1 => lbl4_n_52, B2 => y_address(2), ZN => lbl4_n_78);
  lbl4_g7966 : AOI22D0BWP7T port map(A1 => lbl4_n_63, A2 => lbl4_n_16, B1 => lbl4_n_55, B2 => lbl4_n_20, ZN => lbl4_n_77);
  lbl4_g7967 : OAI22D0BWP7T port map(A1 => lbl4_n_60, A2 => lbl4_n_15, B1 => lbl4_n_57, B2 => lbl4_n_21, ZN => lbl4_n_76);
  lbl4_g7968 : INVD0BWP7T port map(I => lbl4_n_73, ZN => lbl4_n_72);
  lbl4_g7969 : ND2D1BWP7T port map(A1 => lbl4_n_63, A2 => x_address(1), ZN => lbl4_n_70);
  lbl4_g7970 : OR2D1BWP7T port map(A1 => lbl4_n_48, A2 => y_address(2), Z => lbl4_n_75);
  lbl4_g7971 : NR2D1BWP7T port map(A1 => lbl4_n_57, A2 => map_selected(1), ZN => lbl4_n_74);
  lbl4_g7972 : NR2D1BWP7T port map(A1 => lbl4_n_61, A2 => x_address(1), ZN => lbl4_n_73);
  lbl4_g7973 : NR2D1BWP7T port map(A1 => lbl4_n_58, A2 => lbl4_n_2, ZN => lbl4_n_71);
  lbl4_g7974 : AOI22D0BWP7T port map(A1 => lbl4_n_21, A2 => lbl4_n_3, B1 => lbl4_n_6, B2 => x_address(2), ZN => lbl4_n_65);
  lbl4_g7975 : ND3D0BWP7T port map(A1 => start_position_0(3), A2 => lbl4_n_14, A3 => y_address(3), ZN => lbl4_n_69);
  lbl4_g7976 : ND3D0BWP7T port map(A1 => start_position_0(3), A2 => lbl4_n_4, A3 => y_address(4), ZN => lbl4_n_68);
  lbl4_g7977 : OA21D0BWP7T port map(A1 => lbl4_n_17, A2 => lbl4_n_31, B => lbl4_n_60, Z => lbl4_n_67);
  lbl4_g7978 : OR2D1BWP7T port map(A1 => lbl4_n_45, A2 => lbl4_n_13, Z => lbl4_n_66);
  lbl4_g7979 : INVD0BWP7T port map(I => lbl4_n_60, ZN => lbl4_n_59);
  lbl4_g7980 : INVD0BWP7T port map(I => lbl4_n_56, ZN => lbl4_n_55);
  lbl4_g7981 : INVD1BWP7T port map(I => lbl4_n_54, ZN => lbl4_n_53);
  lbl4_g7982 : NR2D0BWP7T port map(A1 => lbl4_n_38, A2 => y_address(3), ZN => lbl4_n_52);
  lbl4_g7983 : IND2D1BWP7T port map(A1 => lbl4_n_38, B1 => lbl4_n_14, ZN => lbl4_n_64);
  lbl4_g7984 : NR2D0BWP7T port map(A1 => lbl4_n_31, A2 => x_address(2), ZN => lbl4_n_63);
  lbl4_g7985 : NR2D0BWP7T port map(A1 => lbl4_n_39, A2 => lbl4_n_4, ZN => lbl4_n_62);
  lbl4_g7986 : ND2D1BWP7T port map(A1 => lbl4_n_23, A2 => x_address(2), ZN => lbl4_n_61);
  lbl4_g7987 : ND2D1BWP7T port map(A1 => lbl4_n_36, A2 => lbl4_n_3, ZN => lbl4_n_60);
  lbl4_g7988 : ND2D1BWP7T port map(A1 => lbl4_n_27, A2 => y_address(4), ZN => lbl4_n_58);
  lbl4_g7989 : OR2D1BWP7T port map(A1 => lbl4_n_31, A2 => lbl4_n_3, Z => lbl4_n_57);
  lbl4_g7990 : ND2D1BWP7T port map(A1 => lbl4_n_36, A2 => x_address(2), ZN => lbl4_n_56);
  lbl4_g7991 : ND2D1BWP7T port map(A1 => lbl4_n_17, A2 => lbl4_n_9, ZN => lbl4_n_54);
  lbl4_g7992 : INVD0BWP7T port map(I => lbl4_n_50, ZN => lbl4_n_51);
  lbl4_g7993 : INVD1BWP7T port map(I => lbl4_n_42, ZN => lbl4_n_41);
  lbl4_g7994 : ND2D1BWP7T port map(A1 => start_position_1(3), A2 => lbl4_n_10, ZN => start_position_0(2));
  lbl4_g7995 : INR2D1BWP7T port map(A1 => lbl4_n_17, B1 => lbl4_n_31, ZN => lbl4_n_50);
  lbl4_g7996 : ND2D1BWP7T port map(A1 => lbl4_n_17, A2 => lbl4_n_36, ZN => lbl4_n_49);
  lbl4_g7997 : OR2D1BWP7T port map(A1 => lbl4_n_24, A2 => lbl4_n_28, Z => lbl4_n_48);
  lbl4_g7998 : MAOI22D0BWP7T port map(A1 => lbl4_n_8, A2 => y_address(1), B1 => lbl4_n_8, B2 => y_address(1), ZN => lbl4_n_47);
  lbl4_g7999 : NR2XD0BWP7T port map(A1 => lbl4_n_22, A2 => lbl4_n_16, ZN => lbl4_n_46);
  lbl4_g8000 : CKAN2D1BWP7T port map(A1 => lbl4_n_37, A2 => lbl4_n_30, Z => lbl4_n_45);
  lbl4_g8001 : NR3D0BWP7T port map(A1 => lbl4_n_6, A2 => lbl4_n_3, A3 => x_address(3), ZN => lbl4_n_44);
  lbl4_g8002 : ND2D1BWP7T port map(A1 => lbl4_n_17, A2 => lbl4_n_32, ZN => lbl4_n_43);
  lbl4_g8003 : ND2D1BWP7T port map(A1 => lbl4_n_12, A2 => lbl4_n_8, ZN => lbl4_n_42);
  lbl4_g8004 : INVD1BWP7T port map(I => lbl4_n_35, ZN => lbl4_n_34);
  lbl4_g8005 : INVD1BWP7T port map(I => lbl4_n_33, ZN => lbl4_n_32);
  lbl4_g8006 : INVD0BWP7T port map(I => lbl4_n_30, ZN => lbl4_n_29);
  lbl4_g8007 : INVD0BWP7T port map(I => lbl4_n_28, ZN => lbl4_n_27);
  lbl4_g8008 : ND2D0BWP7T port map(A1 => map_selected(1), A2 => map_selected(0), ZN => start_position_1(5));
  lbl4_g8009 : CKND2D1BWP7T port map(A1 => y_address(2), A2 => y_address(4), ZN => lbl4_n_39);
  lbl4_g8010 : CKND2D1BWP7T port map(A1 => y_address(1), A2 => y_address(0), ZN => lbl4_n_38);
  lbl4_g8011 : IND2D1BWP7T port map(A1 => y_address(0), B1 => y_address(1), ZN => lbl4_n_37);
  lbl4_g8012 : NR2D1BWP7T port map(A1 => lbl4_n_7, A2 => x_address(3), ZN => lbl4_n_36);
  lbl4_g8013 : ND2D1BWP7T port map(A1 => lbl4_n_4, A2 => map_selected(0), ZN => lbl4_n_35);
  lbl4_g8014 : ND2D1BWP7T port map(A1 => x_address(4), A2 => x_address(3), ZN => lbl4_n_33);
  lbl4_g8015 : ND2D1BWP7T port map(A1 => lbl4_n_7, A2 => x_address(3), ZN => lbl4_n_31);
  lbl4_g8016 : IND2D1BWP7T port map(A1 => y_address(1), B1 => y_address(0), ZN => lbl4_n_30);
  lbl4_g8017 : ND2D1BWP7T port map(A1 => y_address(3), A2 => map_selected(0), ZN => lbl4_n_28);
  lbl4_g8018 : INVD0BWP7T port map(I => lbl4_n_21, ZN => lbl4_n_20);
  lbl4_g8019 : INVD1BWP7T port map(I => lbl4_n_18, ZN => lbl4_n_19);
  lbl4_g8020 : INVD1BWP7T port map(I => lbl4_n_16, ZN => lbl4_n_15);
  lbl4_g8021 : INVD1BWP7T port map(I => lbl4_n_14, ZN => lbl4_n_13);
  lbl4_g8022 : INVD1BWP7T port map(I => start_position_0(3), ZN => lbl4_n_10);
  lbl4_g8023 : ND2D1BWP7T port map(A1 => lbl4_n_2, A2 => map_selected(0), ZN => start_position_1(3));
  lbl4_g8024 : ND2D1BWP7T port map(A1 => lbl4_n_5, A2 => map_selected(1), ZN => lbl4_n_24);
  lbl4_g8025 : NR2XD0BWP7T port map(A1 => x_address(4), A2 => x_address(3), ZN => lbl4_n_23);
  lbl4_g8026 : NR2D1BWP7T port map(A1 => lbl4_n_9, A2 => x_address(1), ZN => lbl4_n_22);
  lbl4_g8027 : ND2D1BWP7T port map(A1 => lbl4_n_6, A2 => lbl4_n_9, ZN => lbl4_n_21);
  lbl4_g8028 : NR2D1BWP7T port map(A1 => lbl4_n_6, A2 => lbl4_n_9, ZN => lbl4_n_18);
  lbl4_g8029 : NR2D1BWP7T port map(A1 => x_address(2), A2 => x_address(1), ZN => lbl4_n_17);
  lbl4_g8030 : NR2D1BWP7T port map(A1 => lbl4_n_6, A2 => x_address(0), ZN => lbl4_n_16);
  lbl4_g8031 : NR2D1BWP7T port map(A1 => lbl4_n_8, A2 => y_address(4), ZN => lbl4_n_14);
  lbl4_g8032 : NR2D1BWP7T port map(A1 => y_address(0), A2 => y_address(1), ZN => lbl4_n_12);
  lbl4_g8033 : NR2XD0BWP7T port map(A1 => lbl4_n_2, A2 => map_selected(0), ZN => start_position_0(3));
  lbl4_g8034 : INVD1BWP7T port map(I => x_address(0), ZN => lbl4_n_9);
  lbl4_g8035 : INVD1BWP7T port map(I => y_address(2), ZN => lbl4_n_8);
  lbl4_g8036 : INVD1BWP7T port map(I => x_address(4), ZN => lbl4_n_7);
  lbl4_g8037 : INVD1BWP7T port map(I => x_address(1), ZN => lbl4_n_6);
  lbl4_g8038 : INVD1BWP7T port map(I => y_address(4), ZN => lbl4_n_5);
  lbl4_g8039 : INVD0BWP7T port map(I => y_address(3), ZN => lbl4_n_4);
  lbl4_g8040 : INVD1BWP7T port map(I => x_address(2), ZN => lbl4_n_3);
  lbl4_g8041 : INVD1BWP7T port map(I => map_selected(1), ZN => lbl4_n_2);
  lbl2_dec1_g100 : AO22D0BWP7T port map(A1 => lbl2_dec1_n_2, A2 => lbl2_data_synced(4), B1 => lbl2_data_synced(5), B2 => lbl2_dec1_n_1, Z => lbl2_walls(6));
  lbl2_dec1_g101 : IOA21D1BWP7T port map(A1 => lbl2_dec1_n_2, A2 => lbl2_dec1_n_0, B => lbl2_dec1_n_5, ZN => lbl2_walls(4));
  lbl2_dec1_g102 : IND2D1BWP7T port map(A1 => lbl2_dec1_n_2, B1 => lbl2_dec1_n_3, ZN => lbl2_walls(5));
  lbl2_dec1_g103 : IOA21D1BWP7T port map(A1 => lbl2_dec1_n_0, A2 => lbl2_data_synced(6), B => lbl2_data_synced(5), ZN => lbl2_dec1_n_5);
  lbl2_dec1_g104 : IOA21D1BWP7T port map(A1 => lbl2_data_synced(6), A2 => lbl2_data_synced(5), B => lbl2_dec1_n_3, ZN => lbl2_walls(7));
  lbl2_dec1_g105 : IND2D1BWP7T port map(A1 => lbl2_data_synced(6), B1 => lbl2_data_synced(4), ZN => lbl2_dec1_n_3);
  lbl2_dec1_g106 : ND2D0BWP7T port map(A1 => lbl2_data_synced(6), A2 => lbl2_data_synced(4), ZN => lbl2_dec1_n_1);
  lbl2_dec1_g107 : INR2D1BWP7T port map(A1 => lbl2_data_synced(6), B1 => lbl2_data_synced(5), ZN => lbl2_dec1_n_2);
  lbl2_dec1_g108 : INVD0BWP7T port map(I => lbl2_data_synced(4), ZN => lbl2_dec1_n_0);
  lbl5_g186 : OAI31D2BWP7T port map(A1 => lbl5_crash_en, A2 => lbl5_engine_en, A3 => lbl5_beep_en, B => FE_OFN5_FE_DBTN24_rst, ZN => lbl5_en0_rst);
  lbl5_g187 : AO31D1BWP7T port map(A1 => pulse_audio, A2 => lbl5_n_2, A3 => lbl5_n_0, B => start_between, Z => lbl5_beep_en);
  lbl5_g188 : AN2D1BWP7T port map(A1 => lbl5_n_2, A2 => game_state(1), Z => lbl5_engine_en);
  lbl5_g189 : IAO21D1BWP7T port map(A1 => game_state(0), A2 => game_state(1), B => game_state(2), ZN => lbl5_crash_en);
  lbl5_g190 : AN2D1BWP7T port map(A1 => game_state(0), A2 => game_state(2), Z => lbl5_n_2);
  lbl5_g192 : INVD0BWP7T port map(I => game_state(1), ZN => lbl5_n_0);
  lbl5_expl_shifter_reg_23 : DFKCNQD1BWP7T port map(CN => FE_PHN46_lbl5_expl_shifter_22, CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => lbl5_expl_shifter(23));
  lbl5_expl_shifter_reg_22 : DFKCNQD1BWP7T port map(CN => FE_PHN59_lbl5_expl_shifter_21, CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => lbl5_expl_shifter(22));
  lbl5_expl_shifter_reg_21 : DFKCNQD1BWP7T port map(CN => FE_PHN49_lbl5_expl_shifter_20, CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => lbl5_expl_shifter(21));
  lbl5_expl_shifter_reg_20 : DFKCNQD1BWP7T port map(CN => FE_PHN33_lbl5_expl_shifter_19, CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => lbl5_expl_shifter(20));
  lbl5_expl_shifter_reg_19 : DFKCNQD1BWP7T port map(CN => lbl5_expl_shifter(18), CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => lbl5_expl_shifter(19));
  lbl5_expl_shifter_reg_18 : DFKCNQD1BWP7T port map(CN => FE_PHN45_lbl5_expl_shifter_17, CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => FE_PHN34_lbl5_expl_shifter_18);
  lbl5_expl_shifter_reg_17 : DFKCNQD1BWP7T port map(CN => FE_PHN44_lbl5_expl_shifter_16, CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => lbl5_expl_shifter(17));
  lbl5_expl_shifter_reg_16 : DFKCNQD1BWP7T port map(CN => lbl5_expl_shifter(15), CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => lbl5_expl_shifter(16));
  lbl5_expl_shifter_reg_15 : DFKCNQD1BWP7T port map(CN => FE_PHN39_lbl5_expl_shifter_14, CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => FE_PHN60_lbl5_expl_shifter_15);
  lbl5_expl_shifter_reg_14 : DFKCNQD1BWP7T port map(CN => FE_PHN41_lbl5_expl_shifter_13, CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => lbl5_expl_shifter(14));
  lbl5_expl_shifter_reg_13 : DFKCNQD1BWP7T port map(CN => lbl5_expl_shifter(12), CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => lbl5_expl_shifter(13));
  lbl5_expl_shifter_reg_12 : DFKCNQD1BWP7T port map(CN => lbl5_expl_shifter(11), CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => FE_PHN37_lbl5_expl_shifter_12);
  lbl5_expl_shifter_reg_11 : DFKCNQD1BWP7T port map(CN => lbl5_expl_shifter(10), CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => FE_PHN40_lbl5_expl_shifter_11);
  lbl5_expl_shifter_reg_10 : DFKCNQD1BWP7T port map(CN => FE_PHN36_lbl5_expl_shifter_9, CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => FE_PHN38_lbl5_expl_shifter_10);
  lbl5_expl_shifter_reg_9 : DFKCNQD1BWP7T port map(CN => FE_PHN35_lbl5_expl_shifter_8, CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => lbl5_expl_shifter(9));
  lbl5_expl_shifter_reg_8 : DFKCNQD1BWP7T port map(CN => lbl5_expl_shifter(7), CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => lbl5_expl_shifter(8));
  lbl5_expl_shifter_reg_7 : DFKCNQD1BWP7T port map(CN => lbl5_expl_shifter(6), CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => FE_PHN43_lbl5_expl_shifter_7);
  lbl5_expl_shifter_reg_6 : DFKCNQD1BWP7T port map(CN => lbl5_expl_shifter(5), CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => FE_PHN58_lbl5_expl_shifter_6);
  lbl5_expl_shifter_reg_5 : DFKCNQD1BWP7T port map(CN => FE_PHN47_lbl5_expl_shifter_4, CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => FE_PHN42_lbl5_expl_shifter_5);
  lbl5_expl_shifter_reg_4 : DFKCNQD1BWP7T port map(CN => lbl5_bits(3), CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => lbl5_expl_shifter(4));
  lbl5_expl_shifter_reg_3 : DFKCNQD1BWP7T port map(CN => lbl5_bits(2), CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => FE_PHN28_lbl5_bits_3);
  lbl5_expl_shifter_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN25_lbl5_bits_1, CP => CTS_21, D => FE_OFN5_FE_DBTN24_rst, Q => FE_PHN27_lbl5_bits_2);
  lbl5_expl_shifter_reg_1 : DFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_19, D => FE_PHN26_lbl5_bits_0, Q => lbl5_bits(1));
  lbl5_expl_shifter_reg_0 : DFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_19, D => FE_PHN295_lbl5_expl_n_1, Q => lbl5_bits(0));
  lbl5_expl_g37 : XNR4D0BWP7T port map(A1 => lbl5_expl_shifter(6), A2 => lbl5_expl_shifter(15), A3 => FE_PHN59_lbl5_expl_shifter_21, A4 => lbl5_expl_shifter(23), ZN => lbl5_expl_n_1);
  lbl5_en0_g2062 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(2), B1 => lbl5_en0_period(3), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_300);
  lbl5_en0_g2063 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => FE_PHN263_lbl5_en0_period_16, B1 => lbl5_en0_period(17), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_314);
  lbl5_en0_g2064 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(14), B1 => lbl5_en0_period(15), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_312);
  lbl5_en0_g2065 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(10), B1 => lbl5_en0_period(11), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_308);
  lbl5_en0_g2066 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(17), B1 => lbl5_en0_period(18), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_315);
  lbl5_en0_g2067 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(9), B1 => lbl5_en0_period(10), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_307);
  lbl5_en0_g2068 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(13), B1 => lbl5_en0_period(14), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_311);
  lbl5_en0_g2069 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(8), B1 => lbl5_en0_period(9), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_306);
  lbl5_en0_g2070 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(5), B1 => lbl5_en0_period(6), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_303);
  lbl5_en0_g2071 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(15), B1 => FE_PHN263_lbl5_en0_period_16, B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_313);
  lbl5_en0_g2072 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(12), B1 => lbl5_en0_period(13), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_310);
  lbl5_en0_g2073 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(6), B1 => lbl5_en0_period(7), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_304);
  lbl5_en0_g2074 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(7), B1 => lbl5_en0_period(8), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_305);
  lbl5_en0_g2075 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(11), B1 => lbl5_en0_period(12), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_309);
  lbl5_en0_g2076 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(4), B1 => lbl5_en0_period(5), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_302);
  lbl5_en0_g2077 : AO22D0BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(3), B1 => lbl5_en0_period(4), B2 => lbl5_en0_frozen_boost, Z => lbl5_en0_n_301);
  lbl5_en0_g2078 : CKAN2D1BWP7T port map(A1 => lbl5_en0_n_278, A2 => lbl5_en0_period(18), Z => lbl5_en0_n_316);
  lbl5_en0_g1824 : MUX2D1BWP7T port map(I0 => lbl5_en0_period(1), I1 => lbl5_en0_period(2), S => lbl5_en0_frozen_boost, Z => lbl5_en0_n_299);
  lbl5_en0_prev_crash_reg : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_crash_en, Q => lbl5_en0_prev_crash);
  lbl5_en0_prev_dir_reg_0 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN171_direction_0_0, Q => lbl5_en0_prev_dir(0));
  lbl5_en0_prev_dir_reg_1 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN255_direction_0_1, Q => lbl5_en0_prev_dir(1));
  lbl5_en0_wave_reg : DFD0BWP7T port map(CP => CTS_19, D => FE_PHN271_lbl5_en0_n_276, Q => UNCONNECTED5, QN => lbl5_en0_n_277);
  lbl5_en0_g3784 : INVD5BWP7T port map(I => lbl5_en0_n_277, ZN => audio(0));
  lbl5_en0_g3785 : OAI211D1BWP7T port map(A1 => lbl5_en0_rst, A2 => lbl5_en0_n_270, B => lbl5_en0_n_327, C => lbl5_en0_n_274, ZN => lbl5_en0_n_276);
  lbl5_en0_g3787 : OAI211D1BWP7T port map(A1 => FE_PHN53_lbl5_en0_frozen_bits_1, A2 => lbl5_en0_n_198, B => lbl5_en0_n_273, C => lbl5_en0_n_269, ZN => lbl5_en0_n_274);
  lbl5_en0_g3788 : AOI211D1BWP7T port map(A1 => lbl5_en0_n_266, A2 => lbl5_en0_count(17), B => lbl5_en0_n_268, C => lbl5_en0_count(18), ZN => lbl5_en0_n_273);
  lbl5_en0_g3789 : IND3D1BWP7T port map(A1 => lbl5_en0_n_280, B1 => lbl5_en0_frozen_bits(3), B2 => lbl5_en0_n_269, ZN => lbl5_en0_n_272);
  lbl5_en0_g3790 : ND3D0BWP7T port map(A1 => lbl5_en0_n_280, A2 => lbl5_en0_n_269, A3 => lbl5_en0_frozen_bits(2), ZN => lbl5_en0_n_271);
  lbl5_en0_g3791 : OAI211D1BWP7T port map(A1 => lbl5_en0_frozen_bits(0), A2 => lbl5_en0_n_198, B => lbl5_en0_n_267, C => lbl5_en0_n_258, ZN => lbl5_en0_n_270);
  lbl5_en0_g3792 : NR3D0BWP7T port map(A1 => lbl5_en0_n_267, A2 => lbl5_en0_rst, A3 => lbl5_en0_n_257, ZN => lbl5_en0_n_269);
  lbl5_en0_g3793 : IAO21D0BWP7T port map(A1 => lbl5_en0_n_266, A2 => lbl5_en0_count(17), B => lbl5_en0_n_316, ZN => lbl5_en0_n_268);
  lbl5_en0_g3794 : NR3D0BWP7T port map(A1 => lbl5_en0_n_265, A2 => lbl5_en0_count(17), A3 => lbl5_en0_count(18), ZN => lbl5_en0_n_267);
  lbl5_en0_g3795 : MAOI222D1BWP7T port map(A => lbl5_en0_n_264, B => lbl5_en0_n_315, C => lbl5_en0_n_196, ZN => lbl5_en0_n_266);
  lbl5_en0_g3796 : MAOI222D1BWP7T port map(A => lbl5_en0_n_263, B => lbl5_en0_n_316, C => lbl5_en0_n_196, ZN => lbl5_en0_n_265);
  lbl5_en0_g3797 : OA221D0BWP7T port map(A1 => lbl5_en0_n_216, A2 => lbl5_en0_n_313, B1 => lbl5_en0_n_191, B2 => lbl5_en0_n_314, C => lbl5_en0_n_261, Z => lbl5_en0_n_264);
  lbl5_en0_g3798 : OA221D0BWP7T port map(A1 => lbl5_en0_n_329, A2 => lbl5_en0_n_314, B1 => lbl5_en0_n_191, B2 => lbl5_en0_n_315, C => lbl5_en0_n_328, Z => lbl5_en0_n_263);
  lbl5_en0_g3800 : AOI32D1BWP7T port map(A1 => lbl5_en0_n_259, A2 => lbl5_en0_n_221, A3 => lbl5_en0_n_204, B1 => lbl5_en0_n_233, B2 => lbl5_en0_n_221, ZN => lbl5_en0_n_261);
  lbl5_en0_g3801 : AOI211XD0BWP7T port map(A1 => lbl5_en0_n_312, A2 => lbl5_en0_n_190, B => lbl5_en0_n_256, C => lbl5_en0_n_207, ZN => lbl5_en0_n_260);
  lbl5_en0_g3802 : AOI32D1BWP7T port map(A1 => lbl5_en0_n_254, A2 => lbl5_en0_n_247, A3 => lbl5_en0_n_234, B1 => lbl5_en0_n_311, B2 => lbl5_en0_n_190, ZN => lbl5_en0_n_259);
  lbl5_en0_g3803 : INVD0BWP7T port map(I => lbl5_en0_n_257, ZN => lbl5_en0_n_258);
  lbl5_en0_g3804 : NR4D0BWP7T port map(A1 => lbl5_en0_n_255, A2 => lbl5_en0_period(17), A3 => lbl5_en0_period(18), A4 => FE_PHN263_lbl5_en0_period_16, ZN => lbl5_en0_n_257);
  lbl5_en0_g3805 : AOI211D1BWP7T port map(A1 => lbl5_en0_n_209, A2 => lbl5_en0_n_199, B => lbl5_en0_n_253, C => lbl5_en0_n_245, ZN => lbl5_en0_n_256);
  lbl5_en0_g3806 : AN3D0BWP7T port map(A1 => lbl5_en0_n_250, A2 => lbl5_en0_period(15), A3 => lbl5_en0_period(14), Z => lbl5_en0_n_255);
  lbl5_en0_g3807 : OAI22D0BWP7T port map(A1 => lbl5_en0_n_251, A2 => lbl5_en0_n_242, B1 => lbl5_en0_n_240, B2 => lbl5_en0_n_237, ZN => lbl5_en0_n_254);
  lbl5_en0_g3808 : AOI31D0BWP7T port map(A1 => lbl5_en0_n_252, A2 => lbl5_en0_n_235, A3 => lbl5_en0_n_222, B => lbl5_en0_n_241, ZN => lbl5_en0_n_253);
  lbl5_en0_g3809 : OA222D0BWP7T port map(A1 => lbl5_en0_n_248, A2 => lbl5_en0_n_225, B1 => lbl5_en0_n_188, B2 => lbl5_en0_n_307, C1 => lbl5_en0_n_304, C2 => lbl5_en0_n_238, Z => lbl5_en0_n_252);
  lbl5_en0_g3810 : OAI222D0BWP7T port map(A1 => lbl5_en0_n_246, A2 => lbl5_en0_n_223, B1 => lbl5_en0_n_303, B2 => lbl5_en0_n_236, C1 => lbl5_en0_n_188, C2 => lbl5_en0_n_306, ZN => lbl5_en0_n_251);
  lbl5_en0_g3811 : AO211D0BWP7T port map(A1 => lbl5_en0_n_249, A2 => lbl5_en0_period(11), B => lbl5_en0_period(13), C => lbl5_en0_period(12), Z => lbl5_en0_n_250);
  lbl5_en0_g3812 : AO211D0BWP7T port map(A1 => lbl5_en0_n_244, A2 => lbl5_en0_period(7), B => lbl5_en0_period(10), C => lbl5_en0_period(9), Z => lbl5_en0_n_249);
  lbl5_en0_g3813 : OAI222D0BWP7T port map(A1 => lbl5_en0_n_231, A2 => lbl5_en0_n_210, B1 => lbl5_en0_count(3), B2 => FE_DBTN12_lbl5_en0_n_303, C1 => lbl5_en0_count(4), C2 => FE_DBTN16_lbl5_en0_n_304, ZN => lbl5_en0_n_248);
  lbl5_en0_g3814 : AOI32D1BWP7T port map(A1 => lbl5_en0_n_214, A2 => FE_DBTN11_lbl5_en0_n_308, A3 => lbl5_en0_count(9), B1 => lbl5_en0_n_240, B2 => lbl5_en0_count(8), ZN => lbl5_en0_n_247);
  lbl5_en0_g3815 : OAI221D0BWP7T port map(A1 => FE_DBTN9_lbl5_en0_n_302, A2 => lbl5_en0_count(3), B1 => lbl5_en0_count(4), B2 => FE_DBTN12_lbl5_en0_n_303, C => lbl5_en0_n_243, ZN => lbl5_en0_n_246);
  lbl5_en0_g3816 : MOAI22D0BWP7T port map(A1 => lbl5_en0_n_226, A2 => lbl5_en0_n_309, B1 => lbl5_en0_n_239, B2 => lbl5_en0_count(8), ZN => lbl5_en0_n_245);
  lbl5_en0_g3817 : OA31D1BWP7T port map(A1 => lbl5_en0_period(6), A2 => lbl5_en0_period(5), A3 => lbl5_en0_n_227, B => lbl5_en0_period(8), Z => lbl5_en0_n_244);
  lbl5_en0_g3818 : AO221D0BWP7T port map(A1 => FE_DBTN17_lbl5_en0_n_301, A2 => lbl5_en0_count(2), B1 => FE_DBTN9_lbl5_en0_n_302, B2 => lbl5_en0_count(3), C => lbl5_en0_n_230, Z => lbl5_en0_n_243);
  lbl5_en0_g3819 : AO33D0BWP7T port map(A1 => lbl5_en0_n_213, A2 => FE_DBTN16_lbl5_en0_n_304, A3 => lbl5_en0_count(5), B1 => lbl5_en0_n_206, B2 => FE_DBTN14_lbl5_en0_n_305, B3 => lbl5_en0_count(6), Z => lbl5_en0_n_242);
  lbl5_en0_g3820 : AOI21D0BWP7T port map(A1 => lbl5_en0_n_224, A2 => lbl5_en0_count(8), B => lbl5_en0_n_239, ZN => lbl5_en0_n_241);
  lbl5_en0_g3821 : IND2D1BWP7T port map(A1 => lbl5_en0_n_225, B1 => lbl5_en0_count(4), ZN => lbl5_en0_n_238);
  lbl5_en0_g3822 : INR2D1BWP7T port map(A1 => lbl5_en0_count(8), B1 => lbl5_en0_n_229, ZN => lbl5_en0_n_237);
  lbl5_en0_g3823 : IND2D1BWP7T port map(A1 => lbl5_en0_n_223, B1 => lbl5_en0_count(4), ZN => lbl5_en0_n_236);
  lbl5_en0_g3824 : NR2D1BWP7T port map(A1 => lbl5_en0_n_229, A2 => lbl5_en0_n_307, ZN => lbl5_en0_n_240);
  lbl5_en0_g3825 : CKAN2D1BWP7T port map(A1 => lbl5_en0_n_224, A2 => FE_DBTN11_lbl5_en0_n_308, Z => lbl5_en0_n_239);
  lbl5_en0_g3826 : ND3D0BWP7T port map(A1 => lbl5_en0_n_220, A2 => FE_DBTN14_lbl5_en0_n_305, A3 => lbl5_en0_count(5), ZN => lbl5_en0_n_235);
  lbl5_en0_g3827 : OAI211D1BWP7T port map(A1 => lbl5_en0_count(11), A2 => lbl5_en0_n_205, B => lbl5_en0_n_208, C => lbl5_en0_n_201, ZN => lbl5_en0_n_234);
  lbl5_en0_g3828 : OAI22D0BWP7T port map(A1 => lbl5_en0_n_215, A2 => lbl5_en0_n_311, B1 => lbl5_en0_n_312, B2 => lbl5_en0_n_193, ZN => lbl5_en0_n_233);
  lbl5_en0_g3829 : OAI32D1BWP7T port map(A1 => lbl5_en0_n_190, A2 => lbl5_en0_n_312, A3 => lbl5_en0_n_207, B1 => lbl5_en0_n_193, B2 => lbl5_en0_n_313, ZN => lbl5_en0_n_232);
  lbl5_en0_g3830 : OA221D0BWP7T port map(A1 => FE_DBTN17_lbl5_en0_n_301, A2 => lbl5_en0_count(1), B1 => lbl5_en0_count(2), B2 => FE_DBTN9_lbl5_en0_n_302, C => lbl5_en0_n_228, Z => lbl5_en0_n_231);
  lbl5_en0_g3831 : OA222D0BWP7T port map(A1 => lbl5_en0_n_218, A2 => lbl5_en0_count(0), B1 => lbl5_en0_count(1), B2 => lbl5_en0_n_186, C1 => lbl5_en0_count(2), C2 => FE_DBTN17_lbl5_en0_n_301, Z => lbl5_en0_n_230);
  lbl5_en0_g3832 : AO211D0BWP7T port map(A1 => FE_DBTN17_lbl5_en0_n_301, A2 => lbl5_en0_count(1), B => lbl5_en0_n_186, C => lbl5_en0_count(0), Z => lbl5_en0_n_228);
  lbl5_en0_g3833 : INR2D1BWP7T port map(A1 => lbl5_en0_period(4), B1 => lbl5_en0_n_211, ZN => lbl5_en0_n_227);
  lbl5_en0_g3834 : ND2D1BWP7T port map(A1 => lbl5_en0_n_219, A2 => lbl5_en0_count(9), ZN => lbl5_en0_n_226);
  lbl5_en0_g3835 : OAI21D0BWP7T port map(A1 => FE_DBTN11_lbl5_en0_n_308, A2 => lbl5_en0_count(9), B => lbl5_en0_n_214, ZN => lbl5_en0_n_229);
  lbl5_en0_g3836 : IND3D1BWP7T port map(A1 => lbl5_en0_n_306, B1 => lbl5_en0_count(6), B2 => lbl5_en0_n_200, ZN => lbl5_en0_n_222);
  lbl5_en0_g3837 : OAI21D0BWP7T port map(A1 => FE_DBTN14_lbl5_en0_n_305, A2 => lbl5_en0_count(5), B => lbl5_en0_n_220, ZN => lbl5_en0_n_225);
  lbl5_en0_g3838 : OA21D0BWP7T port map(A1 => FE_DBTN13_lbl5_en0_n_309, A2 => lbl5_en0_count(9), B => lbl5_en0_n_219, Z => lbl5_en0_n_224);
  lbl5_en0_g3839 : OAI21D0BWP7T port map(A1 => FE_DBTN16_lbl5_en0_n_304, A2 => lbl5_en0_count(5), B => lbl5_en0_n_213, ZN => lbl5_en0_n_223);
  lbl5_en0_g3840 : IOA21D1BWP7T port map(A1 => lbl5_en0_n_186, A2 => lbl5_en0_count(1), B => lbl5_en0_n_299, ZN => lbl5_en0_n_218);
  lbl5_en0_g3842 : ND2D1BWP7T port map(A1 => lbl5_en0_n_202, A2 => lbl5_en0_count(14), ZN => lbl5_en0_n_216);
  lbl5_en0_g3843 : ND2D1BWP7T port map(A1 => lbl5_en0_n_204, A2 => lbl5_en0_count(12), ZN => lbl5_en0_n_215);
  lbl5_en0_g3844 : AOI21D0BWP7T port map(A1 => lbl5_en0_n_313, A2 => lbl5_en0_n_182, B => lbl5_en0_n_203, ZN => lbl5_en0_n_221);
  lbl5_en0_g3845 : OA21D0BWP7T port map(A1 => FE_DBTN15_lbl5_en0_n_306, A2 => lbl5_en0_count(6), B => lbl5_en0_n_200, Z => lbl5_en0_n_220);
  lbl5_en0_g3846 : CKAN2D1BWP7T port map(A1 => lbl5_en0_n_201, A2 => lbl5_en0_n_199, Z => lbl5_en0_n_219);
  lbl5_en0_g3847 : NR4D0BWP7T port map(A1 => lbl5_en0_period(2), A2 => lbl5_en0_period(3), A3 => lbl5_en0_period(1), A4 => lbl5_en0_period(0), ZN => lbl5_en0_n_211);
  lbl5_en0_g3848 : AO22D0BWP7T port map(A1 => FE_DBTN9_lbl5_en0_n_302, A2 => lbl5_en0_count(2), B1 => lbl5_en0_count(3), B2 => FE_DBTN12_lbl5_en0_n_303, Z => lbl5_en0_n_210);
  lbl5_en0_g3849 : AO21D0BWP7T port map(A1 => FE_DBTN10_lbl5_en0_n_311, A2 => lbl5_en0_count(11), B => lbl5_en0_n_205, Z => lbl5_en0_n_209);
  lbl5_en0_g3850 : OAI21D0BWP7T port map(A1 => lbl5_en0_n_310, A2 => lbl5_en0_n_187, B => lbl5_en0_n_309, ZN => lbl5_en0_n_208);
  lbl5_en0_g3851 : MAOI22D0BWP7T port map(A1 => lbl5_en0_n_310, A2 => lbl5_en0_n_187, B1 => FE_DBTN13_lbl5_en0_n_309, B2 => lbl5_en0_count(10), ZN => lbl5_en0_n_214);
  lbl5_en0_g3852 : OA21D0BWP7T port map(A1 => FE_DBTN14_lbl5_en0_n_305, A2 => lbl5_en0_count(6), B => lbl5_en0_n_206, Z => lbl5_en0_n_213);
  lbl5_en0_g3853 : AOI22D0BWP7T port map(A1 => lbl5_en0_n_314, A2 => lbl5_en0_n_182, B1 => lbl5_en0_n_315, B2 => lbl5_en0_n_191, ZN => lbl5_en0_n_212);
  lbl5_en0_g3858 : AN2D1BWP7T port map(A1 => lbl5_en0_n_313, A2 => lbl5_en0_n_193, Z => lbl5_en0_n_207);
  lbl5_en0_g3859 : ND2D1BWP7T port map(A1 => lbl5_en0_n_306, A2 => lbl5_en0_n_188, ZN => lbl5_en0_n_206);
  lbl5_en0_g3860 : INR2XD0BWP7T port map(A1 => lbl5_en0_count(10), B1 => lbl5_en0_n_310, ZN => lbl5_en0_n_205);
  lbl5_en0_g3861 : INVD1BWP7T port map(I => lbl5_en0_n_202, ZN => lbl5_en0_n_203);
  lbl5_en0_g3862 : ND2D1BWP7T port map(A1 => lbl5_en0_n_312, A2 => lbl5_en0_n_193, ZN => lbl5_en0_n_204);
  lbl5_en0_g3863 : ND2D1BWP7T port map(A1 => lbl5_en0_n_314, A2 => lbl5_en0_n_191, ZN => lbl5_en0_n_202);
  lbl5_en0_g3865 : IND2D1BWP7T port map(A1 => lbl5_en0_count(10), B1 => lbl5_en0_n_310, ZN => lbl5_en0_n_201);
  lbl5_en0_g3866 : ND2D1BWP7T port map(A1 => lbl5_en0_n_307, A2 => lbl5_en0_n_188, ZN => lbl5_en0_n_200);
  lbl5_en0_g3867 : ND2D1BWP7T port map(A1 => lbl5_en0_n_311, A2 => lbl5_en0_n_187, ZN => lbl5_en0_n_199);
  lbl5_en0_g3868 : IND2D1BWP7T port map(A1 => lbl5_beep_en, B1 => lbl5_crash_en, ZN => lbl5_en0_n_198);
  lbl5_en0_g3879 : INVD1BWP7T port map(I => lbl5_en0_n_300, ZN => lbl5_en0_n_186);
  lbl5_en0_count_reg_1 : DFKCNQD1BWP7T port map(CN => FE_PHN188_lbl5_en0_n_281, CP => CTS_21, D => lbl5_en0_n_75, Q => lbl5_en0_count(1));
  lbl5_en0_count_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN177_lbl5_en0_n_282, CP => CTS_21, D => lbl5_en0_n_75, Q => lbl5_en0_count(2));
  lbl5_en0_count_reg_3 : DFKCNQD1BWP7T port map(CN => lbl5_en0_n_283, CP => CTS_19, D => lbl5_en0_n_75, Q => lbl5_en0_count(3));
  lbl5_en0_count_reg_4 : DFKCNQD1BWP7T port map(CN => FE_PHN165_lbl5_en0_n_284, CP => CTS_19, D => lbl5_en0_n_75, Q => lbl5_en0_count(4));
  lbl5_en0_count_reg_5 : DFKCNQD1BWP7T port map(CN => FE_PHN184_lbl5_en0_n_285, CP => CTS_19, D => lbl5_en0_n_75, Q => lbl5_en0_count(5));
  lbl5_en0_count_reg_6 : DFKCNQD1BWP7T port map(CN => FE_PHN166_lbl5_en0_n_286, CP => CTS_19, D => lbl5_en0_n_75, Q => lbl5_en0_count(6));
  lbl5_en0_count_reg_8 : DFKCNQD1BWP7T port map(CN => FE_PHN169_lbl5_en0_n_288, CP => CTS_19, D => lbl5_en0_n_75, Q => lbl5_en0_count(8));
  lbl5_en0_count_reg_9 : DFKCNQD1BWP7T port map(CN => FE_PHN180_lbl5_en0_n_289, CP => CTS_19, D => lbl5_en0_n_75, Q => lbl5_en0_count(9));
  lbl5_en0_count_reg_10 : DFKCNQD1BWP7T port map(CN => FE_PHN176_lbl5_en0_n_290, CP => CTS_19, D => lbl5_en0_n_75, Q => lbl5_en0_count(10));
  lbl5_en0_frozen_bits_reg_0 : DFXQD1BWP7T port map(CP => CTS_21, DA => lbl5_en0_frozen_bits(0), DB => FE_PHN26_lbl5_bits_0, Q => FE_PHN57_lbl5_en0_frozen_bits_0, SA => lbl5_en0_n_72);
  lbl5_en0_frozen_bits_reg_1 : DFXQD1BWP7T port map(CP => CTS_19, DA => FE_PHN53_lbl5_en0_frozen_bits_1, DB => FE_PHN25_lbl5_bits_1, Q => lbl5_en0_frozen_bits(1), SA => lbl5_en0_n_72);
  lbl5_en0_frozen_bits_reg_2 : DFXQD1BWP7T port map(CP => CTS_19, DA => lbl5_en0_frozen_bits(2), DB => lbl5_bits(2), Q => FE_PHN121_lbl5_en0_frozen_bits_2, SA => lbl5_en0_n_72);
  lbl5_en0_frozen_bits_reg_3 : DFXQD1BWP7T port map(CP => CTS_19, DA => lbl5_en0_frozen_bits(3), DB => lbl5_bits(3), Q => FE_PHN108_lbl5_en0_frozen_bits_3, SA => lbl5_en0_n_72);
  lbl5_en0_new_period_reg_0 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_151, Q => FE_PHN219_lbl5_en0_new_period_0);
  lbl5_en0_new_period_reg_2 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_158, Q => FE_PHN246_lbl5_en0_new_period_2);
  lbl5_en0_new_period_reg_4 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_168, Q => FE_PHN242_lbl5_en0_new_period_4);
  lbl5_en0_new_period_reg_5 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_169, Q => lbl5_en0_new_period(5));
  lbl5_en0_new_period_reg_6 : DFQD0BWP7T port map(CP => CTS_21, D => lbl5_en0_n_149, Q => FE_PHN341_lbl5_en0_new_period_6);
  lbl5_en0_new_period_reg_8 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_159, Q => lbl5_en0_new_period(8));
  lbl5_en0_new_period_reg_10 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_162, Q => lbl5_en0_new_period(10));
  lbl5_en0_new_period_reg_11 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_166, Q => lbl5_en0_new_period(11));
  lbl5_en0_new_period_reg_14 : DFQD0BWP7T port map(CP => CTS_21, D => lbl5_en0_n_170, Q => FE_PHN243_lbl5_en0_new_period_14);
  lbl5_en0_new_period_reg_15 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_176, Q => FE_PHN202_lbl5_en0_new_period_15);
  lbl5_en0_new_period_reg_16 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_178, Q => FE_PHN192_lbl5_en0_new_period_16);
  lbl5_en0_new_period_reg_18 : DFXQD1BWP7T port map(CP => CTS_21, DA => lbl5_en0_n_177, DB => lbl5_en0_n_174, Q => FE_PHN30_lbl5_en0_new_period_18, SA => lbl5_en0_new_period(18));
  lbl5_en0_period_reg_0 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_98, Q => lbl5_en0_period(0));
  lbl5_en0_period_reg_1 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_92, Q => lbl5_en0_period(1));
  lbl5_en0_period_reg_2 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_91, Q => lbl5_en0_period(2));
  lbl5_en0_period_reg_3 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_90, Q => lbl5_en0_period(3));
  lbl5_en0_period_reg_4 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_80, Q => lbl5_en0_period(4));
  lbl5_en0_period_reg_5 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_89, Q => lbl5_en0_period(5));
  lbl5_en0_period_reg_6 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_88, Q => lbl5_en0_period(6));
  lbl5_en0_period_reg_7 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_87, Q => lbl5_en0_period(7));
  lbl5_en0_period_reg_8 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_95, Q => lbl5_en0_period(8));
  lbl5_en0_period_reg_9 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_86, Q => lbl5_en0_period(9));
  lbl5_en0_period_reg_10 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en0_n_85, Q => lbl5_en0_period(10));
  lbl5_en0_period_reg_11 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_84, Q => lbl5_en0_period(11));
  lbl5_en0_period_reg_12 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en0_n_96, Q => lbl5_en0_period(12));
  lbl5_en0_period_reg_13 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_83, Q => lbl5_en0_period(13));
  lbl5_en0_period_reg_14 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_93, Q => lbl5_en0_period(14));
  lbl5_en0_period_reg_15 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_97, Q => lbl5_en0_period(15));
  lbl5_en0_period_reg_16 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_94, Q => lbl5_en0_period(16));
  lbl5_en0_period_reg_17 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_82, Q => FE_PHN261_lbl5_en0_period_17);
  lbl5_en0_period_reg_18 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_81, Q => FE_PHN264_lbl5_en0_period_18);
  lbl5_en0_g6144 : OAI221D0BWP7T port map(A1 => lbl5_en0_n_175, A2 => FE_PHN111_lbl5_en0_n_8, B1 => FE_PHN64_lbl5_en0_new_period_17, B2 => lbl5_en0_n_173, C => lbl5_en0_n_60, ZN => lbl5_en0_n_179);
  lbl5_en0_g6145 : IND4D0BWP7T port map(A1 => lbl5_en0_n_59, B1 => lbl5_en0_n_3, B2 => lbl5_en0_n_127, B3 => lbl5_en0_n_172, ZN => lbl5_en0_n_178);
  lbl5_en0_g6147 : OAI221D0BWP7T port map(A1 => lbl5_en0_n_109, A2 => FE_PHN64_lbl5_en0_new_period_17, B1 => FE_PHN111_lbl5_en0_n_8, B2 => lbl5_en0_n_111, C => lbl5_en0_n_175, ZN => lbl5_en0_n_177);
  lbl5_en0_g6148 : ND3D0BWP7T port map(A1 => lbl5_en0_n_171, A2 => lbl5_en0_n_163, A3 => lbl5_en0_n_3, ZN => lbl5_en0_n_176);
  lbl5_en0_g6149 : OAI32D1BWP7T port map(A1 => FE_PHN111_lbl5_en0_n_8, A2 => lbl5_en0_n_109, A3 => lbl5_en0_n_160, B1 => FE_PHN64_lbl5_en0_new_period_17, B2 => lbl5_en0_n_127, ZN => lbl5_en0_n_174);
  lbl5_en0_g6150 : AOI221D0BWP7T port map(A1 => lbl5_en0_n_160, A2 => lbl5_en0_n_110, B1 => lbl5_en0_n_112, B2 => lbl5_en0_new_period(16), C => lbl5_en0_n_135, ZN => lbl5_en0_n_175);
  lbl5_en0_g6151 : OA21D0BWP7T port map(A1 => lbl5_en0_n_160, A2 => lbl5_en0_n_109, B => lbl5_en0_n_127, Z => lbl5_en0_n_173);
  lbl5_en0_g6152 : AOI22D0BWP7T port map(A1 => lbl5_en0_n_135, A2 => lbl5_en0_new_period(16), B1 => lbl5_en0_n_167, B2 => lbl5_en0_n_110, ZN => lbl5_en0_n_172);
  lbl5_en0_g6154 : AOI22D0BWP7T port map(A1 => lbl5_en0_n_164, A2 => lbl5_en0_new_period(15), B1 => lbl5_en0_n_59, B2 => FE_PHN171_direction_0_0, ZN => lbl5_en0_n_171);
  lbl5_en0_g6158 : ND3D0BWP7T port map(A1 => lbl5_en0_n_154, A2 => lbl5_en0_n_147, A3 => lbl5_en0_n_3, ZN => lbl5_en0_n_170);
  lbl5_en0_g6162 : AO211D0BWP7T port map(A1 => lbl5_en0_n_145, A2 => FE_PHN318_lbl5_en0_new_period_5, B => lbl5_en0_n_122, C => lbl5_en0_n_115, Z => lbl5_en0_n_169);
  lbl5_en0_g6163 : ND2D1BWP7T port map(A1 => FE_PHN270_lbl5_en0_n_155, A2 => lbl5_en0_n_60, ZN => lbl5_en0_n_168);
  lbl5_en0_g6169 : MOAI22D0BWP7T port map(A1 => lbl5_en0_n_153, A2 => lbl5_en0_new_period(16), B1 => lbl5_en0_n_153, B2 => lbl5_en0_new_period(16), ZN => lbl5_en0_n_167);
  lbl5_en0_g6170 : AO211D0BWP7T port map(A1 => lbl5_en0_n_141, A2 => FE_PHN233_lbl5_en0_new_period_11, B => lbl5_en0_n_116, C => lbl5_en0_n_117, Z => lbl5_en0_n_166);
  lbl5_en0_g6171 : OAI211D1BWP7T port map(A1 => FE_PHN51_lbl5_en0_n_9, A2 => lbl5_en0_n_142, B => lbl5_en0_n_124, C => lbl5_en0_n_60, ZN => lbl5_en0_n_165);
  lbl5_en0_g6172 : AO221D0BWP7T port map(A1 => lbl5_en0_n_119, A2 => lbl5_en0_n_110, B1 => lbl5_en0_n_112, B2 => lbl5_en0_new_period(14), C => lbl5_en0_n_131, Z => lbl5_en0_n_164);
  lbl5_en0_g6173 : AOI22D0BWP7T port map(A1 => lbl5_en0_n_112, A2 => lbl5_en0_n_107, B1 => lbl5_en0_n_152, B2 => lbl5_en0_n_110, ZN => lbl5_en0_n_163);
  lbl5_en0_g6174 : AO221D0BWP7T port map(A1 => lbl5_en0_n_148, A2 => FE_PHN234_lbl5_en0_new_period_10, B1 => lbl5_en0_n_112, B2 => lbl5_en0_n_74, C => lbl5_en0_n_114, Z => lbl5_en0_n_162);
  lbl5_en0_g6175 : OAI211D1BWP7T port map(A1 => FE_PHN52_lbl5_en0_n_14, A2 => lbl5_en0_n_143, B => lbl5_en0_n_123, C => lbl5_en0_n_3, ZN => FE_PHN282_lbl5_en0_n_161);
  lbl5_en0_g6176 : AO211D0BWP7T port map(A1 => lbl5_en0_n_140, A2 => FE_PHN237_lbl5_en0_new_period_8, B => lbl5_en0_n_118, C => lbl5_en0_n_113, Z => lbl5_en0_n_159);
  lbl5_en0_g6177 : IND2D1BWP7T port map(A1 => lbl5_en0_n_153, B1 => lbl5_en0_new_period(16), ZN => lbl5_en0_n_160);
  lbl5_en0_g6181 : MUX2ND0BWP7T port map(I0 => lbl5_en0_n_128, I1 => lbl5_en0_n_144, S => lbl5_en0_new_period(2), ZN => FE_PHN267_lbl5_en0_n_158);
  lbl5_en0_g6182 : OAI21D0BWP7T port map(A1 => lbl5_en0_n_138, A2 => lbl5_en0_n_11, B => lbl5_en0_n_128, ZN => FE_PHN285_lbl5_en0_n_157);
  lbl5_en0_g6183 : OAI211D1BWP7T port map(A1 => FE_PHN118_lbl5_en0_n_6, A2 => lbl5_en0_n_129, B => lbl5_en0_n_136, C => lbl5_en0_n_60, ZN => lbl5_en0_n_156);
  lbl5_en0_g6184 : AOI222D0BWP7T port map(A1 => lbl5_en0_n_139, A2 => lbl5_en0_new_period(4), B1 => lbl5_en0_n_112, B2 => lbl5_en0_n_56, C1 => lbl5_en0_n_110, C2 => lbl5_en0_n_47, ZN => lbl5_en0_n_155);
  lbl5_en0_g6185 : AOI22D0BWP7T port map(A1 => lbl5_en0_n_126, A2 => lbl5_en0_n_110, B1 => lbl5_en0_n_112, B2 => lbl5_en0_n_101, ZN => lbl5_en0_n_154);
  lbl5_en0_g6186 : NR2D1BWP7T port map(A1 => lbl5_en0_n_119, A2 => lbl5_en0_new_period(15), ZN => lbl5_en0_n_152);
  lbl5_en0_g6187 : OAI211D1BWP7T port map(A1 => lbl5_en0_new_period(0), A2 => lbl5_en0_n_111, B => lbl5_en0_n_130, C => lbl5_en0_n_4, ZN => lbl5_en0_n_151);
  lbl5_en0_g6188 : IND2D1BWP7T port map(A1 => lbl5_en0_n_119, B1 => lbl5_en0_new_period(15), ZN => lbl5_en0_n_153);
  lbl5_en0_g6189 : OAI222D0BWP7T port map(A1 => lbl5_en0_n_133, A2 => lbl5_en0_n_7, B1 => FE_PHN292_lbl5_en0_n_46, B2 => lbl5_en0_n_111, C1 => lbl5_en0_n_38, C2 => lbl5_en0_n_120, ZN => lbl5_en0_n_150);
  lbl5_en0_g6190 : AO21D0BWP7T port map(A1 => lbl5_en0_n_132, A2 => FE_PHN265_lbl5_en0_new_period_6, B => lbl5_en0_n_137, Z => lbl5_en0_n_149);
  lbl5_en0_g6191 : AO221D0BWP7T port map(A1 => lbl5_en0_n_110, A2 => lbl5_en0_n_5, B1 => lbl5_en0_n_112, B2 => lbl5_en0_new_period(9), C => lbl5_en0_n_146, Z => lbl5_en0_n_148);
  lbl5_en0_g6192 : AOI22D0BWP7T port map(A1 => lbl5_en0_n_131, A2 => lbl5_en0_new_period(14), B1 => lbl5_en0_n_59, B2 => FE_PHN255_direction_0_1, ZN => lbl5_en0_n_147);
  lbl5_en0_g6193 : OAI221D0BWP7T port map(A1 => lbl5_en0_n_111, A2 => lbl5_en0_n_56, B1 => lbl5_en0_n_0, B2 => lbl5_en0_n_109, C => lbl5_en0_n_104, ZN => lbl5_en0_n_145);
  lbl5_en0_g6194 : AOI221D0BWP7T port map(A1 => lbl5_en0_n_112, A2 => lbl5_en0_n_17, B1 => lbl5_en0_n_110, B2 => lbl5_en0_new_period(1), C => lbl5_en0_n_134, ZN => lbl5_en0_n_144);
  lbl5_en0_g6195 : OA221D0BWP7T port map(A1 => lbl5_en0_n_106, A2 => lbl5_en0_n_109, B1 => FE_PHN118_lbl5_en0_n_6, B2 => lbl5_en0_n_111, C => lbl5_en0_n_129, Z => lbl5_en0_n_143);
  lbl5_en0_g6196 : AOI221D0BWP7T port map(A1 => lbl5_en0_n_110, A2 => lbl5_en0_n_55, B1 => lbl5_en0_n_112, B2 => FE_PHN265_lbl5_en0_new_period_6, C => lbl5_en0_n_132, ZN => lbl5_en0_n_142);
  lbl5_en0_g6197 : AO221D0BWP7T port map(A1 => lbl5_en0_n_112, A2 => lbl5_en0_n_70, B1 => lbl5_en0_n_110, B2 => lbl5_en0_n_69, C => lbl5_en0_n_105, Z => lbl5_en0_n_146);
  lbl5_en0_g6198 : OAI221D0BWP7T port map(A1 => lbl5_en0_n_111, A2 => lbl5_en0_n_74, B1 => lbl5_en0_n_109, B2 => lbl5_en0_n_2, C => lbl5_en0_n_104, ZN => lbl5_en0_n_141);
  lbl5_en0_g6199 : OAI221D0BWP7T port map(A1 => lbl5_en0_n_111, A2 => lbl5_en0_n_64, B1 => lbl5_en0_n_65, B2 => lbl5_en0_n_109, C => lbl5_en0_n_104, ZN => lbl5_en0_n_140);
  lbl5_en0_g6200 : OAI211D1BWP7T port map(A1 => lbl5_en0_n_41, A2 => lbl5_en0_n_111, B => lbl5_en0_n_133, C => lbl5_en0_n_120, ZN => lbl5_en0_n_139);
  lbl5_en0_g6201 : AOI21D0BWP7T port map(A1 => lbl5_en0_n_112, A2 => lbl5_en0_new_period(0), B => lbl5_en0_n_134, ZN => lbl5_en0_n_138);
  lbl5_en0_g6202 : OAI22D0BWP7T port map(A1 => lbl5_en0_n_109, A2 => lbl5_en0_n_57, B1 => lbl5_en0_n_121, B2 => FE_PHN265_lbl5_en0_new_period_6, ZN => lbl5_en0_n_137);
  lbl5_en0_g6203 : AOI22D0BWP7T port map(A1 => lbl5_en0_n_103, A2 => lbl5_en0_n_110, B1 => lbl5_en0_n_117, B2 => FE_PHN118_lbl5_en0_n_6, ZN => lbl5_en0_n_136);
  lbl5_en0_g6204 : OAI21D0BWP7T port map(A1 => lbl5_en0_n_110, A2 => lbl5_en0_n_105, B => lbl5_en0_new_period(0), ZN => lbl5_en0_n_130);
  lbl5_en0_g6205 : OAI21D0BWP7T port map(A1 => lbl5_en0_n_111, A2 => lbl5_en0_n_107, B => lbl5_en0_n_104, ZN => lbl5_en0_n_135);
  lbl5_en0_g6206 : OAI21D0BWP7T port map(A1 => lbl5_en0_n_109, A2 => lbl5_crash_en, B => lbl5_en0_n_104, ZN => lbl5_en0_n_134);
  lbl5_en0_g6207 : AOI21D0BWP7T port map(A1 => lbl5_en0_n_110, A2 => lbl5_en0_n_38, B => lbl5_en0_n_105, ZN => lbl5_en0_n_133);
  lbl5_en0_g6208 : OAI21D0BWP7T port map(A1 => lbl5_en0_n_111, A2 => lbl5_en0_n_61, B => lbl5_en0_n_104, ZN => lbl5_en0_n_132);
  lbl5_en0_g6209 : OAI21D0BWP7T port map(A1 => lbl5_en0_n_111, A2 => lbl5_en0_n_99, B => lbl5_en0_n_104, ZN => lbl5_en0_n_131);
  lbl5_en0_g6210 : MOAI22D0BWP7T port map(A1 => lbl5_en0_n_108, A2 => lbl5_en0_new_period(14), B1 => lbl5_en0_n_108, B2 => lbl5_en0_new_period(14), ZN => lbl5_en0_n_126);
  lbl5_en0_g6211 : OAI22D0BWP7T port map(A1 => lbl5_en0_n_111, A2 => lbl5_en0_n_70, B1 => lbl5_en0_n_109, B2 => lbl5_en0_n_69, ZN => lbl5_en0_n_125);
  lbl5_en0_g6212 : AOI22D0BWP7T port map(A1 => lbl5_en0_n_112, A2 => lbl5_en0_n_64, B1 => lbl5_en0_n_110, B2 => lbl5_en0_n_66, ZN => lbl5_en0_n_124);
  lbl5_en0_g6213 : AOI32D1BWP7T port map(A1 => lbl5_en0_n_106, A2 => lbl5_en0_n_110, A3 => FE_PHN52_lbl5_en0_n_14, B1 => lbl5_en0_n_112, B2 => lbl5_en0_n_99, ZN => lbl5_en0_n_123);
  lbl5_en0_g6214 : AOI21D0BWP7T port map(A1 => lbl5_en0_n_112, A2 => lbl5_en0_n_79, B => lbl5_en0_n_105, ZN => lbl5_en0_n_129);
  lbl5_en0_g6215 : AOI32D1BWP7T port map(A1 => lbl5_en0_n_110, A2 => lbl5_crash_en, A3 => lbl5_en0_n_11, B1 => lbl5_en0_n_112, B2 => lbl5_en0_n_18, ZN => lbl5_en0_n_128);
  lbl5_en0_g6216 : IND3D1BWP7T port map(A1 => lbl5_en0_new_period(16), B1 => lbl5_en0_n_107, B2 => lbl5_en0_n_112, ZN => lbl5_en0_n_127);
  lbl5_en0_g6217 : INVD1BWP7T port map(I => lbl5_en0_n_121, ZN => lbl5_en0_n_122);
  lbl5_en0_g6218 : CKND2D0BWP7T port map(A1 => lbl5_en0_n_112, A2 => lbl5_en0_n_61, ZN => lbl5_en0_n_121);
  lbl5_en0_g6219 : ND2D1BWP7T port map(A1 => lbl5_en0_n_110, A2 => lbl5_en0_n_7, ZN => lbl5_en0_n_120);
  lbl5_en0_g6220 : NR2D0BWP7T port map(A1 => lbl5_en0_n_111, A2 => lbl5_en0_n_70, ZN => lbl5_en0_n_118);
  lbl5_en0_g6221 : IND2D1BWP7T port map(A1 => lbl5_en0_n_108, B1 => lbl5_en0_new_period(14), ZN => lbl5_en0_n_119);
  lbl5_en0_g6222 : INR3D0BWP7T port map(A1 => lbl5_en0_n_2, B1 => FE_PHN233_lbl5_en0_new_period_11, B2 => lbl5_en0_n_109, ZN => lbl5_en0_n_116);
  lbl5_en0_g6223 : INR3D0BWP7T port map(A1 => lbl5_en0_n_0, B1 => FE_PHN249_lbl5_en0_new_period_5, B2 => lbl5_en0_n_109, ZN => lbl5_en0_n_115);
  lbl5_en0_g6224 : NR4D0BWP7T port map(A1 => lbl5_en0_n_109, A2 => lbl5_en0_n_69, A3 => lbl5_en0_n_5, A4 => FE_PHN234_lbl5_en0_new_period_10, ZN => lbl5_en0_n_114);
  lbl5_en0_g6225 : INR3D0BWP7T port map(A1 => lbl5_en0_n_65, B1 => FE_PHN237_lbl5_en0_new_period_8, B2 => lbl5_en0_n_109, ZN => lbl5_en0_n_113);
  lbl5_en0_g6226 : NR2D0BWP7T port map(A1 => lbl5_en0_n_111, A2 => lbl5_en0_n_79, ZN => lbl5_en0_n_117);
  lbl5_en0_g6227 : INVD1BWP7T port map(I => lbl5_en0_n_112, ZN => lbl5_en0_n_111);
  lbl5_en0_g6228 : INVD1BWP7T port map(I => lbl5_en0_n_110, ZN => lbl5_en0_n_109);
  lbl5_en0_g6229 : INR2D1BWP7T port map(A1 => lbl5_engine_en, B1 => lbl5_en0_n_102, ZN => lbl5_en0_n_112);
  lbl5_en0_g6230 : NR2D1BWP7T port map(A1 => lbl5_en0_n_102, A2 => lbl5_engine_en, ZN => lbl5_en0_n_110);
  lbl5_en0_g6231 : ND2D1BWP7T port map(A1 => lbl5_en0_n_106, A2 => FE_PHN236_lbl5_en0_new_period_13, ZN => lbl5_en0_n_108);
  lbl5_en0_g6232 : INR2XD0BWP7T port map(A1 => lbl5_en0_n_101, B1 => lbl5_en0_new_period(15), ZN => lbl5_en0_n_107);
  lbl5_en0_g6233 : INVD1BWP7T port map(I => lbl5_en0_n_105, ZN => lbl5_en0_n_104);
  lbl5_en0_g6234 : HA1D0BWP7T port map(A => lbl5_en0_new_period(12), B => lbl5_en0_n_78, CO => lbl5_en0_n_106, S => lbl5_en0_n_103);
  lbl5_en0_g6236 : NR2D1BWP7T port map(A1 => lbl5_en0_n_62, A2 => lbl5_en0_n_100, ZN => lbl5_en0_n_105);
  lbl5_en0_g6237 : IND2D1BWP7T port map(A1 => lbl5_en0_n_62, B1 => lbl5_en0_n_100, ZN => lbl5_en0_n_102);
  lbl5_en0_g6238 : INR2XD0BWP7T port map(A1 => lbl5_en0_n_99, B1 => lbl5_en0_new_period(14), ZN => lbl5_en0_n_101);
  lbl5_en0_g6249 : AO221D0BWP7T port map(A1 => lbl5_en0_n_77, A2 => lbl5_en0_new_period(0), B1 => lbl5_en0_n_75, B2 => FE_PHN88_lbl5_en0_period_0, C => lbl5_en0_rst, Z => lbl5_en0_n_98);
  lbl5_en0_g6257 : NR4D0BWP7T port map(A1 => lbl5_en0_n_73, A2 => lbl5_en0_count(5), A3 => lbl5_en0_count(6), A4 => lbl5_en0_count(7), ZN => lbl5_en0_n_100);
  lbl5_en0_g6259 : NR3D0BWP7T port map(A1 => lbl5_en0_n_79, A2 => FE_PHN236_lbl5_en0_new_period_13, A3 => lbl5_en0_new_period(12), ZN => lbl5_en0_n_99);
  lbl5_en0_g6281 : AO22D0BWP7T port map(A1 => lbl5_en0_n_77, A2 => lbl5_en0_new_period(15), B1 => FE_PHN91_lbl5_en0_period_15, B2 => lbl5_en0_n_75, Z => lbl5_en0_n_97);
  lbl5_en0_g6282 : MOAI22D0BWP7T port map(A1 => lbl5_en0_n_76, A2 => FE_PHN118_lbl5_en0_n_6, B1 => lbl5_en0_n_75, B2 => FE_PHN105_lbl5_en0_period_12, ZN => lbl5_en0_n_96);
  lbl5_en0_g6283 : AO22D0BWP7T port map(A1 => lbl5_en0_n_77, A2 => FE_PHN237_lbl5_en0_new_period_8, B1 => FE_PHN97_lbl5_en0_period_8, B2 => lbl5_en0_n_75, Z => lbl5_en0_n_95);
  lbl5_en0_g6284 : AO22D0BWP7T port map(A1 => lbl5_en0_n_77, A2 => lbl5_en0_new_period(16), B1 => FE_PHN263_lbl5_en0_period_16, B2 => lbl5_en0_n_75, Z => lbl5_en0_n_94);
  lbl5_en0_g6285 : AO22D0BWP7T port map(A1 => lbl5_en0_n_77, A2 => lbl5_en0_new_period(14), B1 => FE_PHN107_lbl5_en0_period_14, B2 => lbl5_en0_n_75, Z => lbl5_en0_n_93);
  lbl5_en0_g6286 : MOAI22D0BWP7T port map(A1 => lbl5_en0_n_76, A2 => lbl5_en0_n_11, B1 => lbl5_en0_n_75, B2 => FE_PHN63_lbl5_en0_period_1, ZN => lbl5_en0_n_92);
  lbl5_en0_g6287 : AO22D0BWP7T port map(A1 => lbl5_en0_n_77, A2 => lbl5_en0_new_period(2), B1 => FE_PHN98_lbl5_en0_period_2, B2 => lbl5_en0_n_75, Z => lbl5_en0_n_91);
  lbl5_en0_g6288 : MOAI22D0BWP7T port map(A1 => lbl5_en0_n_76, A2 => lbl5_en0_n_7, B1 => lbl5_en0_n_75, B2 => FE_PHN110_lbl5_en0_period_3, ZN => lbl5_en0_n_90);
  lbl5_en0_g6289 : AO22D0BWP7T port map(A1 => lbl5_en0_n_77, A2 => FE_PHN318_lbl5_en0_new_period_5, B1 => FE_PHN124_lbl5_en0_period_5, B2 => lbl5_en0_n_75, Z => lbl5_en0_n_89);
  lbl5_en0_g6290 : AO22D0BWP7T port map(A1 => lbl5_en0_n_77, A2 => FE_PHN265_lbl5_en0_new_period_6, B1 => FE_PHN92_lbl5_en0_period_6, B2 => lbl5_en0_n_75, Z => lbl5_en0_n_88);
  lbl5_en0_g6291 : MOAI22D0BWP7T port map(A1 => lbl5_en0_n_76, A2 => FE_PHN51_lbl5_en0_n_9, B1 => lbl5_en0_n_75, B2 => FE_PHN338_lbl5_en0_period_7, ZN => lbl5_en0_n_87);
  lbl5_en0_g6292 : MOAI22D0BWP7T port map(A1 => lbl5_en0_n_76, A2 => FE_PHN100_lbl5_en0_n_5, B1 => lbl5_en0_n_75, B2 => FE_PHN115_lbl5_en0_period_9, ZN => lbl5_en0_n_86);
  lbl5_en0_g6293 : AO22D0BWP7T port map(A1 => lbl5_en0_n_77, A2 => FE_PHN234_lbl5_en0_new_period_10, B1 => FE_PHN132_lbl5_en0_period_10, B2 => lbl5_en0_n_75, Z => lbl5_en0_n_85);
  lbl5_en0_g6294 : AO22D0BWP7T port map(A1 => lbl5_en0_n_77, A2 => FE_PHN233_lbl5_en0_new_period_11, B1 => FE_PHN72_lbl5_en0_period_11, B2 => lbl5_en0_n_75, Z => lbl5_en0_n_84);
  lbl5_en0_g6295 : MOAI22D0BWP7T port map(A1 => lbl5_en0_n_76, A2 => FE_PHN52_lbl5_en0_n_14, B1 => lbl5_en0_n_75, B2 => FE_PHN144_lbl5_en0_period_13, ZN => lbl5_en0_n_83);
  lbl5_en0_g6296 : MOAI22D0BWP7T port map(A1 => lbl5_en0_n_76, A2 => FE_PHN111_lbl5_en0_n_8, B1 => lbl5_en0_n_75, B2 => lbl5_en0_period(17), ZN => lbl5_en0_n_82);
  lbl5_en0_g6297 : AO22D0BWP7T port map(A1 => lbl5_en0_n_77, A2 => lbl5_en0_new_period(18), B1 => lbl5_en0_period(18), B2 => lbl5_en0_n_75, Z => lbl5_en0_n_81);
  lbl5_en0_g6298 : AO22D0BWP7T port map(A1 => lbl5_en0_n_77, A2 => lbl5_en0_new_period(4), B1 => FE_PHN80_lbl5_en0_period_4, B2 => lbl5_en0_n_75, Z => lbl5_en0_n_80);
  lbl5_en0_g6302 : IND2D1BWP7T port map(A1 => FE_PHN233_lbl5_en0_new_period_11, B1 => lbl5_en0_n_74, ZN => lbl5_en0_n_79);
  lbl5_en0_g6303 : CKAN2D1BWP7T port map(A1 => lbl5_en0_n_2, A2 => FE_PHN233_lbl5_en0_new_period_11, Z => lbl5_en0_n_78);
  lbl5_en0_g6304 : INVD1BWP7T port map(I => lbl5_en0_n_77, ZN => lbl5_en0_n_76);
  lbl5_en0_g6305 : NR2XD0BWP7T port map(A1 => lbl5_en0_n_72, A2 => lbl5_en0_rst, ZN => lbl5_en0_n_77);
  lbl5_en0_g6306 : NR2XD1BWP7T port map(A1 => lbl5_en0_n_71, A2 => lbl5_en0_rst, ZN => lbl5_en0_n_75);
  lbl5_en0_g6307 : IND3D1BWP7T port map(A1 => lbl5_en0_count(4), B1 => lbl5_en0_n_12, B2 => lbl5_en0_n_68, ZN => lbl5_en0_n_73);
  lbl5_en0_g6309 : NR3D0BWP7T port map(A1 => lbl5_en0_n_70, A2 => lbl5_en0_new_period(9), A3 => FE_PHN234_lbl5_en0_new_period_10, ZN => lbl5_en0_n_74);
  lbl5_en0_g6310 : INVD0BWP7T port map(I => lbl5_en0_n_72, ZN => lbl5_en0_n_71);
  lbl5_en0_g6311 : OAI221D1BWP7T port map(A1 => lbl5_en0_n_316, A2 => lbl5_en0_n_10, B1 => lbl5_en0_n_13, B2 => lbl5_en0_n_315, C => lbl5_en0_n_67, ZN => lbl5_en0_n_72);
  lbl5_en0_g6312 : IND2D1BWP7T port map(A1 => FE_PHN237_lbl5_en0_new_period_8, B1 => lbl5_en0_n_64, ZN => lbl5_en0_n_70);
  lbl5_en0_g6313 : ND2D1BWP7T port map(A1 => lbl5_en0_n_65, A2 => FE_PHN237_lbl5_en0_new_period_8, ZN => lbl5_en0_n_69);
  lbl5_en0_g6314 : NR4D0BWP7T port map(A1 => lbl5_en0_n_58, A2 => lbl5_en0_count(3), A3 => lbl5_en0_count(2), A4 => lbl5_en0_count(1), ZN => lbl5_en0_n_68);
  lbl5_en0_g6315 : NR4D0BWP7T port map(A1 => lbl5_en0_n_63, A2 => lbl5_en0_n_42, A3 => lbl5_en0_n_45, A4 => lbl5_en0_n_23, ZN => lbl5_en0_n_67);
  lbl5_en0_g6316 : NR2D0BWP7T port map(A1 => lbl5_en0_n_55, A2 => lbl5_en0_new_period(7), ZN => lbl5_en0_n_66);
  lbl5_en0_g6317 : NR2XD0BWP7T port map(A1 => lbl5_en0_n_55, A2 => lbl5_en0_n_9, ZN => lbl5_en0_n_65);
  lbl5_en0_g6318 : INR3D0BWP7T port map(A1 => lbl5_en0_n_61, B1 => FE_PHN265_lbl5_en0_new_period_6, B2 => lbl5_en0_new_period(7), ZN => lbl5_en0_n_64);
  lbl5_en0_g6319 : ND4D0BWP7T port map(A1 => lbl5_en0_n_53, A2 => lbl5_en0_n_43, A3 => lbl5_en0_n_33, A4 => lbl5_en0_n_36, ZN => lbl5_en0_n_63);
  lbl5_en0_g6320 : ND3D0BWP7T port map(A1 => lbl5_en0_n_4, A2 => lbl5_en0_n_54, A3 => lbl5_en0_n_16, ZN => lbl5_en0_n_62);
  lbl5_en0_g6322 : INR2XD0BWP7T port map(A1 => lbl5_en0_n_56, B1 => FE_PHN249_lbl5_en0_new_period_5, ZN => lbl5_en0_n_61);
  lbl5_en0_g6323 : IND2D1BWP7T port map(A1 => lbl5_en0_n_54, B1 => lbl5_en0_n_4, ZN => lbl5_en0_n_60);
  lbl5_en0_g6324 : OAI21D0BWP7T port map(A1 => lbl5_en0_n_49, A2 => lbl5_en0_frozen_boost, B => lbl5_en0_n_48, ZN => lbl5_en0_n_58);
  lbl5_en0_g6325 : MAOI22D0BWP7T port map(A1 => lbl5_en0_n_51, A2 => lbl5_en0_new_period(6), B1 => lbl5_en0_n_51, B2 => lbl5_en0_new_period(6), ZN => lbl5_en0_n_57);
  lbl5_en0_g6326 : NR3D0BWP7T port map(A1 => lbl5_en0_rst, A2 => lbl5_beep_en, A3 => lbl5_en0_n_52, ZN => lbl5_en0_n_59);
  lbl5_en0_g6327 : INR2XD0BWP7T port map(A1 => lbl5_en0_n_41, B1 => lbl5_en0_new_period(4), ZN => lbl5_en0_n_56);
  lbl5_en0_g6328 : IND2D1BWP7T port map(A1 => lbl5_en0_n_51, B1 => FE_PHN265_lbl5_en0_new_period_6, ZN => lbl5_en0_n_55);
  lbl5_en0_g6329 : AOI21D0BWP7T port map(A1 => lbl5_en0_n_315, A2 => lbl5_en0_n_13, B => lbl5_en0_n_50, ZN => lbl5_en0_n_53);
  lbl5_en0_g6330 : INR2XD0BWP7T port map(A1 => lbl5_en0_n_52, B1 => lbl5_beep_en, ZN => lbl5_en0_n_54);
  lbl5_en0_g6331 : OAI31D0BWP7T port map(A1 => lbl5_en0_n_15, A2 => lbl5_en0_n_19, A3 => lbl5_en0_n_21, B => lbl5_engine_en, ZN => lbl5_en0_n_52);
  lbl5_en0_g6332 : ND2D1BWP7T port map(A1 => lbl5_en0_n_0, A2 => FE_PHN249_lbl5_en0_new_period_5, ZN => lbl5_en0_n_51);
  lbl5_en0_g6333 : OAI211D1BWP7T port map(A1 => lbl5_en0_count(0), A2 => lbl5_en0_n_1, B => lbl5_en0_n_44, C => lbl5_en0_n_24, ZN => lbl5_en0_n_50);
  lbl5_en0_g6334 : AOI31D0BWP7T port map(A1 => lbl5_en0_n_35, A2 => lbl5_en0_n_10, A3 => lbl5_en0_n_13, B => lbl5_en0_count(8), ZN => lbl5_en0_n_49);
  lbl5_en0_g6335 : ND3D0BWP7T port map(A1 => lbl5_en0_n_40, A2 => lbl5_en0_n_13, A3 => lbl5_en0_frozen_boost, ZN => lbl5_en0_n_48);
  lbl5_en0_g6336 : NR3D0BWP7T port map(A1 => lbl5_en0_n_38, A2 => lbl5_en0_n_7, A3 => lbl5_en0_new_period(4), ZN => lbl5_en0_n_47);
  lbl5_en0_g6337 : AOI21D0BWP7T port map(A1 => lbl5_en0_n_39, A2 => lbl5_en0_new_period(3), B => lbl5_en0_n_41, ZN => lbl5_en0_n_46);
  lbl5_en0_g6339 : ND4D0BWP7T port map(A1 => lbl5_en0_n_20, A2 => lbl5_en0_n_30, A3 => lbl5_en0_n_34, A4 => lbl5_en0_n_37, ZN => lbl5_en0_n_45);
  lbl5_en0_g6340 : AOI211XD0BWP7T port map(A1 => lbl5_en0_n_1, A2 => lbl5_en0_count(0), B => lbl5_en0_n_27, C => lbl5_en0_n_28, ZN => lbl5_en0_n_44);
  lbl5_en0_g6341 : AOI211XD0BWP7T port map(A1 => lbl5_en0_n_316, A2 => lbl5_en0_n_10, B => lbl5_en0_n_32, C => lbl5_en0_n_29, ZN => lbl5_en0_n_43);
  lbl5_en0_g6342 : ND4D0BWP7T port map(A1 => lbl5_en0_n_25, A2 => lbl5_en0_n_26, A3 => lbl5_en0_n_22, A4 => lbl5_en0_n_31, ZN => lbl5_en0_n_42);
  lbl5_en0_g6343 : NR2XD0BWP7T port map(A1 => lbl5_en0_n_39, A2 => lbl5_en0_new_period(3), ZN => lbl5_en0_n_41);
  lbl5_en0_g6344 : AOI31D0BWP7T port map(A1 => lbl5_en0_count(13), A2 => lbl5_en0_count(15), A3 => lbl5_en0_count(14), B => lbl5_en0_count(16), ZN => lbl5_en0_n_40);
  lbl5_en0_g6345 : XNR2D1BWP7T port map(A1 => lbl5_en0_n_313, A2 => lbl5_en0_count(15), ZN => lbl5_en0_n_37);
  lbl5_en0_g6346 : XNR2D1BWP7T port map(A1 => lbl5_en0_n_305, A2 => lbl5_en0_count(7), ZN => lbl5_en0_n_36);
  lbl5_en0_g6347 : ND3D0BWP7T port map(A1 => lbl5_en0_count(15), A2 => lbl5_en0_count(16), A3 => lbl5_en0_count(14), ZN => lbl5_en0_n_35);
  lbl5_en0_g6348 : XNR2D1BWP7T port map(A1 => lbl5_en0_n_312, A2 => lbl5_en0_count(14), ZN => lbl5_en0_n_34);
  lbl5_en0_g6349 : XNR2D1BWP7T port map(A1 => lbl5_en0_n_302, A2 => lbl5_en0_count(4), ZN => lbl5_en0_n_33);
  lbl5_en0_g6350 : CKXOR2D1BWP7T port map(A1 => lbl5_en0_n_303, A2 => lbl5_en0_count(5), Z => lbl5_en0_n_32);
  lbl5_en0_g6351 : XNR2D1BWP7T port map(A1 => lbl5_en0_n_309, A2 => lbl5_en0_count(11), ZN => lbl5_en0_n_31);
  lbl5_en0_g6352 : XNR2D1BWP7T port map(A1 => lbl5_en0_n_310, A2 => lbl5_en0_count(12), ZN => lbl5_en0_n_30);
  lbl5_en0_g6353 : IND2D1BWP7T port map(A1 => lbl5_en0_new_period(2), B1 => lbl5_en0_n_18, ZN => lbl5_en0_n_39);
  lbl5_en0_g6355 : OAI21D0BWP7T port map(A1 => lbl5_en0_new_period(2), A2 => lbl5_en0_new_period(1), B => lbl5_crash_en, ZN => lbl5_en0_n_38);
  lbl5_en0_g6356 : CKXOR2D1BWP7T port map(A1 => lbl5_en0_n_304, A2 => lbl5_en0_count(6), Z => lbl5_en0_n_29);
  lbl5_en0_g6357 : CKXOR2D1BWP7T port map(A1 => lbl5_en0_n_299, A2 => lbl5_en0_count(1), Z => lbl5_en0_n_28);
  lbl5_en0_g6358 : CKXOR2D1BWP7T port map(A1 => lbl5_en0_n_300, A2 => lbl5_en0_count(2), Z => lbl5_en0_n_27);
  lbl5_en0_g6359 : XNR2D1BWP7T port map(A1 => lbl5_en0_n_307, A2 => lbl5_en0_count(9), ZN => lbl5_en0_n_26);
  lbl5_en0_g6360 : XNR2D1BWP7T port map(A1 => lbl5_en0_n_306, A2 => lbl5_en0_count(8), ZN => lbl5_en0_n_25);
  lbl5_en0_g6361 : XNR2D1BWP7T port map(A1 => lbl5_en0_n_301, A2 => lbl5_en0_count(3), ZN => lbl5_en0_n_24);
  lbl5_en0_g6362 : CKXOR2D1BWP7T port map(A1 => lbl5_en0_n_314, A2 => lbl5_en0_count(16), Z => lbl5_en0_n_23);
  lbl5_en0_g6363 : XNR2D1BWP7T port map(A1 => lbl5_en0_n_308, A2 => lbl5_en0_count(10), ZN => lbl5_en0_n_22);
  lbl5_en0_g6364 : CKXOR2D1BWP7T port map(A1 => FE_PHN255_direction_0_1, A2 => lbl5_en0_prev_dir(1), Z => lbl5_en0_n_21);
  lbl5_en0_g6365 : XNR2D1BWP7T port map(A1 => lbl5_en0_n_311, A2 => lbl5_en0_count(13), ZN => lbl5_en0_n_20);
  lbl5_en0_g6366 : CKXOR2D1BWP7T port map(A1 => direction_0(0), A2 => lbl5_en0_prev_dir(0), Z => lbl5_en0_n_19);
  lbl5_en0_g6367 : INVD0BWP7T port map(I => lbl5_en0_n_18, ZN => lbl5_en0_n_17);
  lbl5_en0_g6368 : NR2XD0BWP7T port map(A1 => lbl5_en0_new_period(0), A2 => lbl5_en0_new_period(1), ZN => lbl5_en0_n_18);
  lbl5_en0_g6370 : IND2D1BWP7T port map(A1 => lbl5_en0_prev_crash, B1 => lbl5_crash_en, ZN => lbl5_en0_n_16);
  lbl5_en0_g6385 : INVD1BWP7T port map(I => lbl5_en0_rst, ZN => lbl5_en0_n_4);
  lbl5_en0_g2 : IND3D1BWP7T port map(A1 => FE_PHN56_lbl5_en0_n_16, B1 => lbl5_en0_n_4, B2 => lbl5_en0_n_54, ZN => lbl5_en0_n_3);
  lbl5_en0_g6386 : INR3D0BWP7T port map(A1 => FE_PHN234_lbl5_en0_new_period_10, B1 => lbl5_en0_n_69, B2 => lbl5_en0_n_5, ZN => lbl5_en0_n_2);
  lbl5_en0_g6387 : MUX2ND0BWP7T port map(I0 => lbl5_en0_period(0), I1 => lbl5_en0_period(1), S => lbl5_en0_frozen_boost, ZN => lbl5_en0_n_1);
  lbl5_en0_g6388 : INR3D0BWP7T port map(A1 => lbl5_en0_new_period(4), B1 => lbl5_en0_n_38, B2 => lbl5_en0_n_7, ZN => lbl5_en0_n_0);
  lbl5_en0_g6389 : AO211D0BWP7T port map(A1 => lbl5_en0_n_272, A2 => lbl5_en0_n_271, B => lbl5_en0_n_198, C => lbl5_en0_n_273, Z => lbl5_en0_n_327);
  lbl5_en0_g6390 : OAI21D0BWP7T port map(A1 => lbl5_en0_n_232, A2 => lbl5_en0_n_260, B => lbl5_en0_n_212, ZN => lbl5_en0_n_328);
  lbl5_en0_frozen_boost_reg : DFXD1BWP7T port map(CP => CTS_19, DA => FE_PHN199_lbl5_en0_frozen_boost, DB => FE_PHN104_boost_audio_0, Q => lbl5_en0_frozen_boost, QN => lbl5_en0_n_278, SA => lbl5_en0_n_72);
  lbl5_en0_count_reg_16 : DFKCND1BWP7T port map(CN => lbl5_en0_n_75, CP => CTS_19, D => lbl5_en0_n_296, Q => FE_PHN254_lbl5_en0_count_16, QN => lbl5_en0_n_196);
  lbl5_en0_count_reg_13 : DFKCND1BWP7T port map(CN => lbl5_en0_n_293, CP => CTS_19, D => lbl5_en0_n_75, Q => lbl5_en0_count(13), QN => lbl5_en0_n_193);
  lbl5_en0_count_reg_15 : DFKCND1BWP7T port map(CN => lbl5_en0_n_75, CP => CTS_19, D => FE_PHN141_lbl5_en0_n_295, Q => lbl5_en0_count(15), QN => lbl5_en0_n_191);
  lbl5_en0_count_reg_12 : DFKCND1BWP7T port map(CN => lbl5_en0_n_292, CP => CTS_19, D => lbl5_en0_n_75, Q => lbl5_en0_count(12), QN => lbl5_en0_n_190);
  lbl5_en0_count_reg_7 : DFKCND1BWP7T port map(CN => lbl5_en0_n_287, CP => CTS_19, D => lbl5_en0_n_75, Q => lbl5_en0_count(7), QN => lbl5_en0_n_188);
  lbl5_en0_count_reg_11 : DFKCND1BWP7T port map(CN => FE_PHN175_lbl5_en0_n_291, CP => CTS_19, D => lbl5_en0_n_75, Q => lbl5_en0_count(11), QN => lbl5_en0_n_187);
  lbl5_en0_count_reg_14 : DFKCND1BWP7T port map(CN => lbl5_en0_n_75, CP => CTS_19, D => FE_PHN158_lbl5_en0_n_294, Q => lbl5_en0_count(14), QN => lbl5_en0_n_182);
  lbl5_en0_prev_engine_reg : DFD1BWP7T port map(CP => CTS_21, D => lbl5_engine_en, Q => lbl5_en0_prev_engine, QN => lbl5_en0_n_15);
  lbl5_en0_new_period_reg_13 : DFD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_161, Q => lbl5_en0_new_period(13), QN => lbl5_en0_n_14);
  lbl5_en0_count_reg_17 : DFKCND1BWP7T port map(CN => lbl5_en0_n_75, CP => CTS_19, D => lbl5_en0_n_297, Q => FE_PHN251_lbl5_en0_count_17, QN => lbl5_en0_n_13);
  lbl5_en0_count_reg_0 : DFKCND1BWP7T port map(CN => FE_PHN62_lbl5_en0_n_12, CP => CTS_19, D => lbl5_en0_n_75, Q => lbl5_en0_count(0), QN => lbl5_en0_n_12);
  lbl5_en0_new_period_reg_1 : DFD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_157, Q => lbl5_en0_new_period(1), QN => FE_PHN54_lbl5_en0_n_11);
  lbl5_en0_count_reg_18 : DFKCND1BWP7T port map(CN => lbl5_en0_n_75, CP => CTS_19, D => FE_PHN281_lbl5_en0_n_298, Q => lbl5_en0_count(18), QN => lbl5_en0_n_10);
  lbl5_en0_new_period_reg_7 : DFD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_165, Q => FE_PHN220_lbl5_en0_new_period_7, QN => lbl5_en0_n_9);
  lbl5_en0_new_period_reg_17 : DFD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_179, Q => lbl5_en0_new_period(17), QN => lbl5_en0_n_8);
  lbl5_en0_new_period_reg_3 : DFD1BWP7T port map(CP => CTS_21, D => lbl5_en0_n_150, Q => lbl5_en0_new_period(3), QN => FE_PHN329_lbl5_en0_n_7);
  lbl5_en0_new_period_reg_12 : DFD1BWP7T port map(CP => CTS_21, D => FE_PHN284_lbl5_en0_n_156, Q => lbl5_en0_new_period(12), QN => lbl5_en0_n_6);
  lbl5_en0_new_period_reg_9 : DFXD1BWP7T port map(CP => CTS_21, DA => lbl5_en0_n_146, DB => lbl5_en0_n_125, Q => FE_PHN230_lbl5_en0_new_period_9, QN => lbl5_en0_n_5, SA => lbl5_en0_new_period(9));
  lbl5_en0_g6429 : IOA21D0BWP7T port map(A1 => lbl5_en0_n_315, A2 => lbl5_en0_n_191, B => lbl5_en0_count(14), ZN => lbl5_en0_n_329);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1075 : AN4D1BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_34, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_31, A3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_30, A4 => lbl5_en0_csa_tree_lt_140_15_groupi_n_28, Z => lbl5_en0_n_280);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1076 : AOI31D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_27, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_37, A3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_54, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_33, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_34);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1077 : ND4D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_32, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_24, A3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_21, A4 => lbl5_en0_csa_tree_lt_140_15_groupi_n_23, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_33);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1078 : IND3D0BWP7T port map(A1 => lbl5_en0_n_301, B1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_36, B2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_29, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_32);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1079 : OAI211D1BWP7T port map(A1 => FE_DBTN17_lbl5_en0_n_301, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_36, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_29, C => lbl5_en0_csa_tree_lt_140_15_groupi_n_4, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_31);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1080 : AOI33D1BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_26, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_38, A3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_55, B1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_20, B2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_41, B3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_58, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_30);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1081 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_37, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_54, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_27, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_29);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1082 : AOI33D1BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_25, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_39, A3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_56, B1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_22, B2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_40, B3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_57, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_28);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1083 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_38, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_55, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_26, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_27);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1084 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_39, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_56, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_25, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_26);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1085 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_40, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_57, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_22, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_25);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1086 : AOI33D1BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_18, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_42, A3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_59, B1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_13, B2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_45, B3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_62, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_24);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1087 : AOI31D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_8, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_49, A3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_66, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_19, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_23);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1088 : AOI33D1BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_16, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_43, A3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_60, B1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_12, B2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_46, B3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_63, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_21);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1089 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_41, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_58, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_20, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_22);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1090 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_42, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_59, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_18, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_20);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1091 : ND4D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_17, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_14, A3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_10, A4 => lbl5_en0_csa_tree_lt_140_15_groupi_n_6, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_19);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1092 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_43, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_60, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_16, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_18);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1093 : ND3D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_15, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_44, A3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_61, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_17);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1094 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_44, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_61, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_15, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_16);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1095 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_45, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_62, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_13, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_15);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1096 : AOI33D1BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_11, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_47, A3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_64, B1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_9, B2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_48, B3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_65, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_14);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1097 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_46, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_63, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_12, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_13);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1098 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_47, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_64, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_11, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_12);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1099 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_48, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_65, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_9, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_11);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1100 : AOI33D1BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_7, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_50, A3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_67, B1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_5, B2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_51, B3 => lbl5_en0_csa_tree_lt_140_15_groupi_n_68, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_10);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1101 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_49, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_66, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_8, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_9);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1102 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_50, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_67, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_7, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_8);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1103 : OA21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_51, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_68, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_5, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_7);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1104 : AOI22D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_3, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_52, B1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_53, B2 => lbl5_en0_count(18), ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_6);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1105 : AO21D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_2, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_52, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_3, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_5);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1106 : MAOI222D1BWP7T port map(A => lbl5_en0_n_300, B => lbl5_en0_n_299, C => lbl5_en0_csa_tree_lt_140_15_groupi_n_0, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_4);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1107 : AN2D0BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_2, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_69, Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_3);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1108 : OR2D1BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_53, A2 => lbl5_en0_count(18), Z => lbl5_en0_csa_tree_lt_140_15_groupi_n_2);
  lbl5_en0_csa_tree_lt_140_15_groupi_g1110 : CKND1BWP7T port map(I => lbl5_en0_count(0), ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_0);
  lbl5_en0_csa_tree_lt_140_15_groupi_g882 : FA1D0BWP7T port map(A => lbl5_en0_csa_tree_lt_140_15_groupi_n_124, B => lbl5_en0_count(16), CI => lbl5_en0_csa_tree_lt_140_15_groupi_n_112, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_69, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_51);
  lbl5_en0_csa_tree_lt_140_15_groupi_g883 : FA1D0BWP7T port map(A => lbl5_en0_csa_tree_lt_140_15_groupi_n_112, B => lbl5_en0_count(15), CI => lbl5_en0_csa_tree_lt_140_15_groupi_n_123, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_68, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_50);
  lbl5_en0_csa_tree_lt_140_15_groupi_g884 : FA1D0BWP7T port map(A => lbl5_en0_csa_tree_lt_140_15_groupi_n_121, B => lbl5_en0_count(13), CI => lbl5_en0_csa_tree_lt_140_15_groupi_n_119, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_66, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_48);
  lbl5_en0_csa_tree_lt_140_15_groupi_g885 : FA1D0BWP7T port map(A => FE_DBTN9_lbl5_en0_n_302, B => lbl5_en0_count(2), CI => FE_DBTN17_lbl5_en0_n_301, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_55, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_37);
  lbl5_en0_csa_tree_lt_140_15_groupi_g886 : FA1D0BWP7T port map(A => FE_DBTN12_lbl5_en0_n_303, B => lbl5_en0_count(3), CI => FE_DBTN9_lbl5_en0_n_302, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_56, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_38);
  lbl5_en0_csa_tree_lt_140_15_groupi_g887 : FA1D0BWP7T port map(A => FE_DBTN16_lbl5_en0_n_304, B => lbl5_en0_count(4), CI => FE_DBTN12_lbl5_en0_n_303, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_57, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_39);
  lbl5_en0_csa_tree_lt_140_15_groupi_g888 : FA1D0BWP7T port map(A => FE_DBTN14_lbl5_en0_n_305, B => lbl5_en0_count(5), CI => FE_DBTN16_lbl5_en0_n_304, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_58, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_40);
  lbl5_en0_csa_tree_lt_140_15_groupi_g889 : FA1D0BWP7T port map(A => FE_DBTN15_lbl5_en0_n_306, B => lbl5_en0_count(6), CI => FE_DBTN14_lbl5_en0_n_305, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_59, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_41);
  lbl5_en0_csa_tree_lt_140_15_groupi_g890 : FA1D0BWP7T port map(A => lbl5_en0_csa_tree_lt_140_15_groupi_n_118, B => lbl5_en0_count(7), CI => FE_DBTN15_lbl5_en0_n_306, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_60, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_42);
  lbl5_en0_csa_tree_lt_140_15_groupi_g891 : FA1D0BWP7T port map(A => FE_DBTN13_lbl5_en0_n_309, B => lbl5_en0_count(9), CI => FE_DBTN11_lbl5_en0_n_308, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_62, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_44);
  lbl5_en0_csa_tree_lt_140_15_groupi_g892 : FA1D0BWP7T port map(A => FE_DBTN11_lbl5_en0_n_308, B => lbl5_en0_count(8), CI => lbl5_en0_csa_tree_lt_140_15_groupi_n_118, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_61, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_43);
  lbl5_en0_csa_tree_lt_140_15_groupi_g893 : FA1D0BWP7T port map(A => lbl5_en0_csa_tree_lt_140_15_groupi_n_120, B => lbl5_en0_count(10), CI => FE_DBTN13_lbl5_en0_n_309, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_63, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_45);
  lbl5_en0_csa_tree_lt_140_15_groupi_g894 : FA1D0BWP7T port map(A => FE_DBTN10_lbl5_en0_n_311, B => lbl5_en0_count(11), CI => lbl5_en0_csa_tree_lt_140_15_groupi_n_120, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_64, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_46);
  lbl5_en0_csa_tree_lt_140_15_groupi_g895 : FA1D0BWP7T port map(A => lbl5_en0_csa_tree_lt_140_15_groupi_n_119, B => lbl5_en0_count(12), CI => FE_DBTN10_lbl5_en0_n_311, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_65, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_47);
  lbl5_en0_csa_tree_lt_140_15_groupi_g896 : FA1D0BWP7T port map(A => lbl5_en0_csa_tree_lt_140_15_groupi_n_123, B => lbl5_en0_count(14), CI => lbl5_en0_csa_tree_lt_140_15_groupi_n_121, CO => lbl5_en0_csa_tree_lt_140_15_groupi_n_67, S => lbl5_en0_csa_tree_lt_140_15_groupi_n_49);
  lbl5_en0_csa_tree_lt_140_15_groupi_g897 : OAI21D0BWP7T port map(A1 => lbl5_en0_n_300, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_114, B => lbl5_en0_csa_tree_lt_140_15_groupi_n_54, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_36);
  lbl5_en0_csa_tree_lt_140_15_groupi_g898 : IOA21D1BWP7T port map(A1 => lbl5_en0_csa_tree_lt_140_15_groupi_n_124, A2 => lbl5_en0_count(17), B => lbl5_en0_csa_tree_lt_140_15_groupi_n_53, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_52);
  lbl5_en0_csa_tree_lt_140_15_groupi_g899 : ND2D1BWP7T port map(A1 => lbl5_en0_n_300, A2 => lbl5_en0_csa_tree_lt_140_15_groupi_n_114, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_54);
  lbl5_en0_csa_tree_lt_140_15_groupi_g900 : IND2D1BWP7T port map(A1 => lbl5_en0_count(17), B1 => lbl5_en0_n_316, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_53);
  lbl5_en0_csa_tree_lt_140_15_groupi_g901 : INVD1BWP7T port map(I => lbl5_en0_n_316, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_124);
  lbl5_en0_csa_tree_lt_140_15_groupi_g902 : INVD0BWP7T port map(I => lbl5_en0_n_314, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_123);
  lbl5_en0_csa_tree_lt_140_15_groupi_g904 : INVD1BWP7T port map(I => lbl5_en0_n_313, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_121);
  lbl5_en0_csa_tree_lt_140_15_groupi_g905 : INVD1BWP7T port map(I => lbl5_en0_n_310, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_120);
  lbl5_en0_csa_tree_lt_140_15_groupi_g906 : INVD1BWP7T port map(I => lbl5_en0_n_312, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_119);
  lbl5_en0_csa_tree_lt_140_15_groupi_g907 : INVD1BWP7T port map(I => lbl5_en0_n_307, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_118);
  lbl5_en0_csa_tree_lt_140_15_groupi_g911 : CKND1BWP7T port map(I => lbl5_en0_count(1), ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_114);
  lbl5_en0_csa_tree_lt_140_15_groupi_g913 : INVD1BWP7T port map(I => lbl5_en0_n_315, ZN => lbl5_en0_csa_tree_lt_140_15_groupi_n_112);
  lbl5_en1_g2069 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(2), B1 => lbl5_en1_period(3), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_304);
  lbl5_en1_g2070 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => FE_PHN259_lbl5_en1_period_16, B1 => lbl5_en1_period(17), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_318);
  lbl5_en1_g2071 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(14), B1 => lbl5_en1_period(15), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_316);
  lbl5_en1_g2072 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(10), B1 => lbl5_en1_period(11), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_312);
  lbl5_en1_g2073 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(17), B1 => lbl5_en1_period(18), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_319);
  lbl5_en1_g2074 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(9), B1 => lbl5_en1_period(10), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_311);
  lbl5_en1_g2075 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(13), B1 => lbl5_en1_period(14), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_315);
  lbl5_en1_g2076 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(8), B1 => lbl5_en1_period(9), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_310);
  lbl5_en1_g2077 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(5), B1 => lbl5_en1_period(6), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_307);
  lbl5_en1_g2078 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(15), B1 => FE_PHN259_lbl5_en1_period_16, B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_317);
  lbl5_en1_g2079 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(12), B1 => lbl5_en1_period(13), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_314);
  lbl5_en1_g2080 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(6), B1 => lbl5_en1_period(7), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_308);
  lbl5_en1_g2081 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(7), B1 => lbl5_en1_period(8), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_309);
  lbl5_en1_g2082 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(11), B1 => lbl5_en1_period(12), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_313);
  lbl5_en1_g2083 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(4), B1 => lbl5_en1_period(5), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_306);
  lbl5_en1_g2084 : AO22D0BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(3), B1 => lbl5_en1_period(4), B2 => lbl5_en1_frozen_boost, Z => lbl5_en1_n_305);
  lbl5_en1_g2085 : CKAN2D1BWP7T port map(A1 => lbl5_en1_n_282, A2 => lbl5_en1_period(18), Z => lbl5_en1_n_320);
  lbl5_en1_g1831 : MUX2D1BWP7T port map(I0 => lbl5_en1_period(1), I1 => lbl5_en1_period(2), S => lbl5_en1_frozen_boost, Z => lbl5_en1_n_303);
  lbl5_en1_prev_crash_reg : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_crash_en, Q => lbl5_en1_prev_crash);
  lbl5_en1_prev_dir_reg_0 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN126_direction_1_0, Q => lbl5_en1_prev_dir(0));
  lbl5_en1_prev_dir_reg_1 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN128_direction_1_1, Q => lbl5_en1_prev_dir(1));
  lbl5_en1_prev_engine_reg : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_engine_en, Q => lbl5_en1_prev_engine);
  lbl5_en1_wave_reg : DFD0BWP7T port map(CP => CTS_19, D => FE_PHN273_lbl5_en1_n_280, Q => UNCONNECTED6, QN => lbl5_en1_n_281);
  lbl5_en1_g3791 : INVD5BWP7T port map(I => lbl5_en1_n_281, ZN => audio(1));
  lbl5_en1_g3792 : OAI211D1BWP7T port map(A1 => lbl5_en0_rst, A2 => lbl5_en1_n_274, B => lbl5_en1_n_331, C => lbl5_en1_n_278, ZN => lbl5_en1_n_280);
  lbl5_en1_g3794 : OAI211D1BWP7T port map(A1 => lbl5_en1_frozen_bits(1), A2 => lbl5_en1_n_202, B => lbl5_en1_n_277, C => lbl5_en1_n_273, ZN => lbl5_en1_n_278);
  lbl5_en1_g3795 : AOI211D1BWP7T port map(A1 => lbl5_en1_n_270, A2 => FE_PHN185_lbl5_en1_count_17, B => lbl5_en1_n_272, C => lbl5_en1_count(18), ZN => lbl5_en1_n_277);
  lbl5_en1_g3796 : IND3D1BWP7T port map(A1 => lbl5_en1_n_284, B1 => lbl5_en1_frozen_bits(3), B2 => lbl5_en1_n_273, ZN => lbl5_en1_n_276);
  lbl5_en1_g3797 : ND3D0BWP7T port map(A1 => lbl5_en1_n_284, A2 => lbl5_en1_n_273, A3 => FE_PHN81_lbl5_en1_frozen_bits_2, ZN => lbl5_en1_n_275);
  lbl5_en1_g3798 : OAI211D1BWP7T port map(A1 => FE_PHN131_lbl5_en1_frozen_bits_0, A2 => lbl5_en1_n_202, B => lbl5_en1_n_271, C => lbl5_en1_n_262, ZN => lbl5_en1_n_274);
  lbl5_en1_g3799 : NR3D0BWP7T port map(A1 => lbl5_en1_n_271, A2 => lbl5_en0_rst, A3 => lbl5_en1_n_261, ZN => lbl5_en1_n_273);
  lbl5_en1_g3800 : IAO21D0BWP7T port map(A1 => lbl5_en1_n_270, A2 => FE_PHN185_lbl5_en1_count_17, B => lbl5_en1_n_320, ZN => lbl5_en1_n_272);
  lbl5_en1_g3801 : NR3D0BWP7T port map(A1 => lbl5_en1_n_269, A2 => FE_PHN185_lbl5_en1_count_17, A3 => lbl5_en1_count(18), ZN => lbl5_en1_n_271);
  lbl5_en1_g3802 : MAOI222D1BWP7T port map(A => lbl5_en1_n_268, B => lbl5_en1_n_319, C => lbl5_en1_n_200, ZN => lbl5_en1_n_270);
  lbl5_en1_g3803 : MAOI222D1BWP7T port map(A => lbl5_en1_n_267, B => lbl5_en1_n_320, C => lbl5_en1_n_200, ZN => lbl5_en1_n_269);
  lbl5_en1_g3804 : OA221D0BWP7T port map(A1 => lbl5_en1_n_220, A2 => lbl5_en1_n_317, B1 => lbl5_en1_n_195, B2 => lbl5_en1_n_318, C => lbl5_en1_n_265, Z => lbl5_en1_n_268);
  lbl5_en1_g3805 : OA221D0BWP7T port map(A1 => lbl5_en1_n_333, A2 => lbl5_en1_n_318, B1 => lbl5_en1_n_195, B2 => lbl5_en1_n_319, C => lbl5_en1_n_332, Z => lbl5_en1_n_267);
  lbl5_en1_g3807 : AOI32D1BWP7T port map(A1 => lbl5_en1_n_263, A2 => lbl5_en1_n_225, A3 => lbl5_en1_n_208, B1 => lbl5_en1_n_237, B2 => lbl5_en1_n_225, ZN => lbl5_en1_n_265);
  lbl5_en1_g3808 : AOI211XD0BWP7T port map(A1 => lbl5_en1_n_316, A2 => lbl5_en1_n_194, B => lbl5_en1_n_260, C => lbl5_en1_n_211, ZN => lbl5_en1_n_264);
  lbl5_en1_g3809 : AOI32D1BWP7T port map(A1 => lbl5_en1_n_258, A2 => lbl5_en1_n_251, A3 => lbl5_en1_n_238, B1 => lbl5_en1_n_315, B2 => lbl5_en1_n_194, ZN => lbl5_en1_n_263);
  lbl5_en1_g3810 : INVD0BWP7T port map(I => lbl5_en1_n_261, ZN => lbl5_en1_n_262);
  lbl5_en1_g3811 : NR4D0BWP7T port map(A1 => lbl5_en1_n_259, A2 => lbl5_en1_period(17), A3 => lbl5_en1_period(18), A4 => FE_PHN259_lbl5_en1_period_16, ZN => lbl5_en1_n_261);
  lbl5_en1_g3812 : AOI211D1BWP7T port map(A1 => lbl5_en1_n_213, A2 => lbl5_en1_n_203, B => lbl5_en1_n_257, C => lbl5_en1_n_249, ZN => lbl5_en1_n_260);
  lbl5_en1_g3813 : AN3D0BWP7T port map(A1 => lbl5_en1_n_254, A2 => lbl5_en1_period(15), A3 => lbl5_en1_period(14), Z => lbl5_en1_n_259);
  lbl5_en1_g3814 : OAI22D0BWP7T port map(A1 => lbl5_en1_n_255, A2 => lbl5_en1_n_246, B1 => lbl5_en1_n_244, B2 => lbl5_en1_n_241, ZN => lbl5_en1_n_258);
  lbl5_en1_g3815 : AOI31D0BWP7T port map(A1 => lbl5_en1_n_256, A2 => lbl5_en1_n_239, A3 => lbl5_en1_n_226, B => lbl5_en1_n_245, ZN => lbl5_en1_n_257);
  lbl5_en1_g3816 : OA222D0BWP7T port map(A1 => lbl5_en1_n_252, A2 => lbl5_en1_n_229, B1 => lbl5_en1_n_192, B2 => lbl5_en1_n_311, C1 => lbl5_en1_n_308, C2 => lbl5_en1_n_242, Z => lbl5_en1_n_256);
  lbl5_en1_g3817 : OAI222D0BWP7T port map(A1 => lbl5_en1_n_250, A2 => lbl5_en1_n_227, B1 => lbl5_en1_n_307, B2 => lbl5_en1_n_240, C1 => lbl5_en1_n_192, C2 => lbl5_en1_n_310, ZN => lbl5_en1_n_255);
  lbl5_en1_g3818 : AO211D0BWP7T port map(A1 => lbl5_en1_n_253, A2 => lbl5_en1_period(11), B => lbl5_en1_period(13), C => lbl5_en1_period(12), Z => lbl5_en1_n_254);
  lbl5_en1_g3819 : AO211D0BWP7T port map(A1 => lbl5_en1_n_248, A2 => lbl5_en1_period(7), B => lbl5_en1_period(10), C => lbl5_en1_period(9), Z => lbl5_en1_n_253);
  lbl5_en1_g3820 : OAI222D0BWP7T port map(A1 => lbl5_en1_n_235, A2 => lbl5_en1_n_214, B1 => lbl5_en1_count(3), B2 => FE_DBTN3_lbl5_en1_n_307, C1 => lbl5_en1_count(4), C2 => FE_DBTN7_lbl5_en1_n_308, ZN => lbl5_en1_n_252);
  lbl5_en1_g3821 : AOI32D1BWP7T port map(A1 => lbl5_en1_n_218, A2 => FE_DBTN2_lbl5_en1_n_312, A3 => lbl5_en1_count(9), B1 => lbl5_en1_n_244, B2 => lbl5_en1_count(8), ZN => lbl5_en1_n_251);
  lbl5_en1_g3822 : OAI221D0BWP7T port map(A1 => FE_DBTN0_lbl5_en1_n_306, A2 => lbl5_en1_count(3), B1 => lbl5_en1_count(4), B2 => FE_DBTN3_lbl5_en1_n_307, C => lbl5_en1_n_247, ZN => lbl5_en1_n_250);
  lbl5_en1_g3823 : MOAI22D0BWP7T port map(A1 => lbl5_en1_n_230, A2 => lbl5_en1_n_313, B1 => lbl5_en1_n_243, B2 => lbl5_en1_count(8), ZN => lbl5_en1_n_249);
  lbl5_en1_g3824 : OA31D1BWP7T port map(A1 => lbl5_en1_period(6), A2 => lbl5_en1_period(5), A3 => lbl5_en1_n_231, B => lbl5_en1_period(8), Z => lbl5_en1_n_248);
  lbl5_en1_g3825 : AO221D0BWP7T port map(A1 => FE_DBTN8_lbl5_en1_n_305, A2 => lbl5_en1_count(2), B1 => FE_DBTN0_lbl5_en1_n_306, B2 => lbl5_en1_count(3), C => lbl5_en1_n_234, Z => lbl5_en1_n_247);
  lbl5_en1_g3826 : AO33D0BWP7T port map(A1 => lbl5_en1_n_217, A2 => FE_DBTN7_lbl5_en1_n_308, A3 => lbl5_en1_count(5), B1 => lbl5_en1_n_210, B2 => FE_DBTN5_lbl5_en1_n_309, B3 => lbl5_en1_count(6), Z => lbl5_en1_n_246);
  lbl5_en1_g3827 : AOI21D0BWP7T port map(A1 => lbl5_en1_n_228, A2 => lbl5_en1_count(8), B => lbl5_en1_n_243, ZN => lbl5_en1_n_245);
  lbl5_en1_g3828 : IND2D1BWP7T port map(A1 => lbl5_en1_n_229, B1 => lbl5_en1_count(4), ZN => lbl5_en1_n_242);
  lbl5_en1_g3829 : INR2D1BWP7T port map(A1 => lbl5_en1_count(8), B1 => lbl5_en1_n_233, ZN => lbl5_en1_n_241);
  lbl5_en1_g3830 : IND2D1BWP7T port map(A1 => lbl5_en1_n_227, B1 => lbl5_en1_count(4), ZN => lbl5_en1_n_240);
  lbl5_en1_g3831 : NR2D1BWP7T port map(A1 => lbl5_en1_n_233, A2 => lbl5_en1_n_311, ZN => lbl5_en1_n_244);
  lbl5_en1_g3832 : CKAN2D1BWP7T port map(A1 => lbl5_en1_n_228, A2 => FE_DBTN2_lbl5_en1_n_312, Z => lbl5_en1_n_243);
  lbl5_en1_g3833 : ND3D0BWP7T port map(A1 => lbl5_en1_n_224, A2 => FE_DBTN5_lbl5_en1_n_309, A3 => lbl5_en1_count(5), ZN => lbl5_en1_n_239);
  lbl5_en1_g3834 : OAI211D1BWP7T port map(A1 => lbl5_en1_count(11), A2 => lbl5_en1_n_209, B => lbl5_en1_n_212, C => lbl5_en1_n_205, ZN => lbl5_en1_n_238);
  lbl5_en1_g3835 : OAI22D0BWP7T port map(A1 => lbl5_en1_n_219, A2 => lbl5_en1_n_315, B1 => lbl5_en1_n_316, B2 => lbl5_en1_n_197, ZN => lbl5_en1_n_237);
  lbl5_en1_g3836 : OAI32D1BWP7T port map(A1 => lbl5_en1_n_194, A2 => lbl5_en1_n_316, A3 => lbl5_en1_n_211, B1 => lbl5_en1_n_197, B2 => lbl5_en1_n_317, ZN => lbl5_en1_n_236);
  lbl5_en1_g3837 : OA221D0BWP7T port map(A1 => FE_DBTN8_lbl5_en1_n_305, A2 => lbl5_en1_count(1), B1 => lbl5_en1_count(2), B2 => FE_DBTN0_lbl5_en1_n_306, C => lbl5_en1_n_232, Z => lbl5_en1_n_235);
  lbl5_en1_g3838 : OA222D0BWP7T port map(A1 => lbl5_en1_n_222, A2 => lbl5_en1_count(0), B1 => lbl5_en1_count(1), B2 => lbl5_en1_n_190, C1 => lbl5_en1_count(2), C2 => FE_DBTN8_lbl5_en1_n_305, Z => lbl5_en1_n_234);
  lbl5_en1_g3839 : AO211D0BWP7T port map(A1 => FE_DBTN8_lbl5_en1_n_305, A2 => lbl5_en1_count(1), B => lbl5_en1_n_190, C => lbl5_en1_count(0), Z => lbl5_en1_n_232);
  lbl5_en1_g3840 : INR2D1BWP7T port map(A1 => lbl5_en1_period(4), B1 => lbl5_en1_n_215, ZN => lbl5_en1_n_231);
  lbl5_en1_g3841 : ND2D1BWP7T port map(A1 => lbl5_en1_n_223, A2 => lbl5_en1_count(9), ZN => lbl5_en1_n_230);
  lbl5_en1_g3842 : OAI21D0BWP7T port map(A1 => FE_DBTN2_lbl5_en1_n_312, A2 => lbl5_en1_count(9), B => lbl5_en1_n_218, ZN => lbl5_en1_n_233);
  lbl5_en1_g3843 : IND3D1BWP7T port map(A1 => lbl5_en1_n_310, B1 => lbl5_en1_count(6), B2 => lbl5_en1_n_204, ZN => lbl5_en1_n_226);
  lbl5_en1_g3844 : OAI21D0BWP7T port map(A1 => FE_DBTN5_lbl5_en1_n_309, A2 => lbl5_en1_count(5), B => lbl5_en1_n_224, ZN => lbl5_en1_n_229);
  lbl5_en1_g3845 : OA21D0BWP7T port map(A1 => FE_DBTN4_lbl5_en1_n_313, A2 => lbl5_en1_count(9), B => lbl5_en1_n_223, Z => lbl5_en1_n_228);
  lbl5_en1_g3846 : OAI21D0BWP7T port map(A1 => FE_DBTN7_lbl5_en1_n_308, A2 => lbl5_en1_count(5), B => lbl5_en1_n_217, ZN => lbl5_en1_n_227);
  lbl5_en1_g3847 : IOA21D1BWP7T port map(A1 => lbl5_en1_n_190, A2 => lbl5_en1_count(1), B => lbl5_en1_n_303, ZN => lbl5_en1_n_222);
  lbl5_en1_g3849 : ND2D1BWP7T port map(A1 => lbl5_en1_n_206, A2 => lbl5_en1_count(14), ZN => lbl5_en1_n_220);
  lbl5_en1_g3850 : ND2D1BWP7T port map(A1 => lbl5_en1_n_208, A2 => lbl5_en1_count(12), ZN => lbl5_en1_n_219);
  lbl5_en1_g3851 : AOI21D0BWP7T port map(A1 => lbl5_en1_n_317, A2 => lbl5_en1_n_186, B => lbl5_en1_n_207, ZN => lbl5_en1_n_225);
  lbl5_en1_g3852 : OA21D0BWP7T port map(A1 => FE_DBTN6_lbl5_en1_n_310, A2 => lbl5_en1_count(6), B => lbl5_en1_n_204, Z => lbl5_en1_n_224);
  lbl5_en1_g3853 : CKAN2D1BWP7T port map(A1 => lbl5_en1_n_205, A2 => lbl5_en1_n_203, Z => lbl5_en1_n_223);
  lbl5_en1_g3854 : NR4D0BWP7T port map(A1 => lbl5_en1_period(2), A2 => lbl5_en1_period(3), A3 => lbl5_en1_period(1), A4 => lbl5_en1_period(0), ZN => lbl5_en1_n_215);
  lbl5_en1_g3855 : AO22D0BWP7T port map(A1 => FE_DBTN0_lbl5_en1_n_306, A2 => lbl5_en1_count(2), B1 => lbl5_en1_count(3), B2 => FE_DBTN3_lbl5_en1_n_307, Z => lbl5_en1_n_214);
  lbl5_en1_g3856 : AO21D0BWP7T port map(A1 => FE_DBTN1_lbl5_en1_n_315, A2 => lbl5_en1_count(11), B => lbl5_en1_n_209, Z => lbl5_en1_n_213);
  lbl5_en1_g3857 : OAI21D0BWP7T port map(A1 => lbl5_en1_n_314, A2 => lbl5_en1_n_191, B => lbl5_en1_n_313, ZN => lbl5_en1_n_212);
  lbl5_en1_g3858 : MAOI22D0BWP7T port map(A1 => lbl5_en1_n_314, A2 => lbl5_en1_n_191, B1 => FE_DBTN4_lbl5_en1_n_313, B2 => lbl5_en1_count(10), ZN => lbl5_en1_n_218);
  lbl5_en1_g3859 : OA21D0BWP7T port map(A1 => FE_DBTN5_lbl5_en1_n_309, A2 => lbl5_en1_count(6), B => lbl5_en1_n_210, Z => lbl5_en1_n_217);
  lbl5_en1_g3860 : AOI22D0BWP7T port map(A1 => lbl5_en1_n_318, A2 => lbl5_en1_n_186, B1 => lbl5_en1_n_319, B2 => lbl5_en1_n_195, ZN => lbl5_en1_n_216);
  lbl5_en1_g3865 : AN2D1BWP7T port map(A1 => lbl5_en1_n_317, A2 => lbl5_en1_n_197, Z => lbl5_en1_n_211);
  lbl5_en1_g3866 : ND2D1BWP7T port map(A1 => lbl5_en1_n_310, A2 => lbl5_en1_n_192, ZN => lbl5_en1_n_210);
  lbl5_en1_g3867 : INR2XD0BWP7T port map(A1 => lbl5_en1_count(10), B1 => lbl5_en1_n_314, ZN => lbl5_en1_n_209);
  lbl5_en1_g3868 : INVD1BWP7T port map(I => lbl5_en1_n_206, ZN => lbl5_en1_n_207);
  lbl5_en1_g3869 : ND2D1BWP7T port map(A1 => lbl5_en1_n_316, A2 => lbl5_en1_n_197, ZN => lbl5_en1_n_208);
  lbl5_en1_g3870 : ND2D1BWP7T port map(A1 => lbl5_en1_n_318, A2 => lbl5_en1_n_195, ZN => lbl5_en1_n_206);
  lbl5_en1_g3872 : IND2D1BWP7T port map(A1 => lbl5_en1_count(10), B1 => lbl5_en1_n_314, ZN => lbl5_en1_n_205);
  lbl5_en1_g3873 : ND2D1BWP7T port map(A1 => lbl5_en1_n_311, A2 => lbl5_en1_n_192, ZN => lbl5_en1_n_204);
  lbl5_en1_g3874 : ND2D1BWP7T port map(A1 => lbl5_en1_n_315, A2 => lbl5_en1_n_191, ZN => lbl5_en1_n_203);
  lbl5_en1_g3875 : IND2D1BWP7T port map(A1 => lbl5_beep_en, B1 => lbl5_crash_en, ZN => lbl5_en1_n_202);
  lbl5_en1_g3886 : INVD1BWP7T port map(I => lbl5_en1_n_304, ZN => lbl5_en1_n_190);
  lbl5_en1_count_reg_1 : DFKCNQD1BWP7T port map(CN => lbl5_en1_n_285, CP => CTS_19, D => lbl5_en1_n_74, Q => lbl5_en1_count(1));
  lbl5_en1_count_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN130_lbl5_en1_n_286, CP => CTS_19, D => lbl5_en1_n_74, Q => lbl5_en1_count(2));
  lbl5_en1_count_reg_3 : DFKCNQD1BWP7T port map(CN => FE_PHN179_lbl5_en1_n_287, CP => CTS_19, D => lbl5_en1_n_74, Q => lbl5_en1_count(3));
  lbl5_en1_count_reg_4 : DFKCNQD1BWP7T port map(CN => FE_PHN183_lbl5_en1_n_288, CP => CTS_19, D => lbl5_en1_n_74, Q => lbl5_en1_count(4));
  lbl5_en1_count_reg_5 : DFKCNQD1BWP7T port map(CN => FE_PHN178_lbl5_en1_n_289, CP => CTS_19, D => lbl5_en1_n_74, Q => lbl5_en1_count(5));
  lbl5_en1_count_reg_6 : DFKCNQD1BWP7T port map(CN => FE_PHN195_lbl5_en1_n_290, CP => CTS_19, D => lbl5_en1_n_74, Q => lbl5_en1_count(6));
  lbl5_en1_count_reg_8 : DFKCNQD1BWP7T port map(CN => FE_PHN189_lbl5_en1_n_292, CP => CTS_19, D => lbl5_en1_n_74, Q => lbl5_en1_count(8));
  lbl5_en1_count_reg_9 : DFKCNQD1BWP7T port map(CN => FE_PHN173_lbl5_en1_n_293, CP => CTS_19, D => lbl5_en1_n_74, Q => lbl5_en1_count(9));
  lbl5_en1_count_reg_10 : DFKCNQD1BWP7T port map(CN => FE_PHN161_lbl5_en1_n_294, CP => CTS_19, D => lbl5_en1_n_74, Q => lbl5_en1_count(10));
  lbl5_en1_frozen_bits_reg_0 : DFXQD1BWP7T port map(CP => CTS_19, DA => FE_PHN26_lbl5_bits_0, DB => FE_PHN131_lbl5_en1_frozen_bits_0, Q => lbl5_en1_frozen_bits(0), SA => lbl5_en1_n_73);
  lbl5_en1_frozen_bits_reg_1 : DFXQD1BWP7T port map(CP => CTS_19, DA => FE_PHN25_lbl5_bits_1, DB => FE_PHN313_lbl5_en1_frozen_bits_1, Q => FE_PHN125_lbl5_en1_frozen_bits_1, SA => lbl5_en1_n_73);
  lbl5_en1_frozen_bits_reg_2 : DFXQD1BWP7T port map(CP => CTS_19, DA => lbl5_bits(2), DB => FE_PHN81_lbl5_en1_frozen_bits_2, Q => lbl5_en1_frozen_bits(2), SA => lbl5_en1_n_73);
  lbl5_en1_frozen_bits_reg_3 : DFXQD1BWP7T port map(CP => CTS_19, DA => lbl5_bits(3), DB => lbl5_en1_frozen_bits(3), Q => FE_PHN96_lbl5_en1_frozen_bits_3, SA => lbl5_en1_n_73);
  lbl5_en1_new_period_reg_1 : DFXQD1BWP7T port map(CP => CTS_19, DA => lbl5_en1_n_144, DB => lbl5_en1_n_133, Q => FE_PHN252_lbl5_en1_new_period_1, SA => FE_PHN321_lbl5_en1_new_period_1);
  lbl5_en1_new_period_reg_2 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_170, Q => lbl5_en1_new_period(2));
  lbl5_en1_new_period_reg_3 : DFQD1BWP7T port map(CP => CTS_20, D => lbl5_en1_n_173, Q => FE_PHN248_lbl5_en1_new_period_3);
  lbl5_en1_new_period_reg_13 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en1_n_178, Q => lbl5_en1_new_period(13));
  lbl5_en1_new_period_reg_14 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN289_lbl5_en1_n_179, Q => lbl5_en1_new_period(14));
  lbl5_en1_new_period_reg_15 : DFQD1BWP7T port map(CP => CTS_21, D => lbl5_en1_n_174, Q => lbl5_en1_new_period(15));
  lbl5_en1_new_period_reg_16 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN287_lbl5_en1_n_183, Q => lbl5_en1_new_period(16));
  lbl5_en1_new_period_reg_18 : DFXQD1BWP7T port map(CP => CTS_19, DA => lbl5_en1_n_171, DB => lbl5_en1_n_1, Q => FE_PHN31_lbl5_en1_new_period_18, SA => lbl5_en1_new_period(18));
  lbl5_en1_period_reg_0 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_100, Q => lbl5_en1_period(0));
  lbl5_en1_period_reg_1 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_93, Q => lbl5_en1_period(1));
  lbl5_en1_period_reg_2 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_92, Q => lbl5_en1_period(2));
  lbl5_en1_period_reg_3 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_91, Q => lbl5_en1_period(3));
  lbl5_en1_period_reg_4 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_90, Q => lbl5_en1_period(4));
  lbl5_en1_period_reg_5 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_89, Q => lbl5_en1_period(5));
  lbl5_en1_period_reg_6 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_83, Q => lbl5_en1_period(6));
  lbl5_en1_period_reg_7 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_88, Q => lbl5_en1_period(7));
  lbl5_en1_period_reg_8 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_81, Q => lbl5_en1_period(8));
  lbl5_en1_period_reg_9 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_80, Q => lbl5_en1_period(9));
  lbl5_en1_period_reg_10 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_94, Q => lbl5_en1_period(10));
  lbl5_en1_period_reg_11 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_87, Q => lbl5_en1_period(11));
  lbl5_en1_period_reg_12 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_97, Q => lbl5_en1_period(12));
  lbl5_en1_period_reg_13 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_96, Q => lbl5_en1_period(13));
  lbl5_en1_period_reg_14 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_85, Q => lbl5_en1_period(14));
  lbl5_en1_period_reg_15 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_84, Q => lbl5_en1_period(15));
  lbl5_en1_period_reg_16 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_82, Q => lbl5_en1_period(16));
  lbl5_en1_period_reg_17 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_86, Q => FE_PHN260_lbl5_en1_period_17);
  lbl5_en1_period_reg_18 : DFQD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_95, Q => lbl5_en1_period(18));
  lbl5_en1_g6864 : IND4D0BWP7T port map(A1 => lbl5_en1_n_65, B1 => lbl5_en1_n_59, B2 => lbl5_en1_n_145, B3 => lbl5_en1_n_172, ZN => lbl5_en1_n_183);
  lbl5_en1_g6875 : ND4D0BWP7T port map(A1 => lbl5_en1_n_164, A2 => lbl5_en1_n_137, A3 => lbl5_en1_n_125, A4 => lbl5_en1_n_59, ZN => FE_PHN278_lbl5_en1_n_182);
  lbl5_en1_g6876 : ND3D0BWP7T port map(A1 => lbl5_en1_n_169, A2 => lbl5_en1_n_124, A3 => lbl5_en1_n_64, ZN => lbl5_en1_n_181);
  lbl5_en1_g6877 : AO211D0BWP7T port map(A1 => lbl5_en1_n_165, A2 => lbl5_en1_new_period(17), B => lbl5_en1_n_162, C => lbl5_en1_n_63, Z => lbl5_en1_n_180);
  lbl5_en1_g6878 : IND3D1BWP7T port map(A1 => lbl5_en1_n_65, B1 => lbl5_en1_n_130, B2 => lbl5_en1_n_167, ZN => lbl5_en1_n_179);
  lbl5_en1_g6880 : OR3D1BWP7T port map(A1 => lbl5_en1_n_65, A2 => lbl5_en1_n_113, A3 => lbl5_en1_n_163, Z => FE_PHN306_lbl5_en1_n_178);
  lbl5_en1_g6881 : OAI211D1BWP7T port map(A1 => lbl5_en1_n_7, A2 => lbl5_en1_n_159, B => lbl5_en1_n_148, C => lbl5_en1_n_64, ZN => lbl5_en1_n_177);
  lbl5_en1_g6884 : OAI211D1BWP7T port map(A1 => lbl5_en1_n_6, A2 => lbl5_en1_n_152, B => lbl5_en1_n_138, C => lbl5_en1_n_114, ZN => lbl5_en1_n_176);
  lbl5_en1_g6885 : OAI211D1BWP7T port map(A1 => FE_PHN223_lbl5_en1_n_8, A2 => lbl5_en1_n_156, B => lbl5_en1_n_135, C => lbl5_en1_n_116, ZN => lbl5_en1_n_175);
  lbl5_en1_g6886 : AO211D0BWP7T port map(A1 => lbl5_en1_n_153, A2 => FE_PHN203_lbl5_en1_new_period_15, B => lbl5_en1_n_160, C => lbl5_en1_n_65, Z => lbl5_en1_n_174);
  lbl5_en1_g6887 : AO211D0BWP7T port map(A1 => lbl5_en1_n_118, A2 => lbl5_en1_n_42, B => lbl5_en1_n_166, C => lbl5_en1_n_143, Z => lbl5_en1_n_173);
  lbl5_en1_g6888 : AOI222D0BWP7T port map(A1 => lbl5_en1_n_161, A2 => FE_PHN213_lbl5_en1_new_period_16, B1 => lbl5_en1_n_129, B2 => FE_PHN203_lbl5_en1_new_period_15, C1 => lbl5_en1_n_105, C2 => lbl5_en1_n_21, ZN => lbl5_en1_n_172);
  lbl5_en1_g6889 : AO221D0BWP7T port map(A1 => lbl5_en1_n_105, A2 => lbl5_en1_new_period(17), B1 => lbl5_en1_n_107, B2 => FE_PHN146_lbl5_en1_n_5, C => lbl5_en1_n_165, Z => lbl5_en1_n_171);
  lbl5_en1_g6894 : AO22D0BWP7T port map(A1 => lbl5_en1_n_157, A2 => FE_PHN244_lbl5_en1_new_period_2, B1 => lbl5_en1_n_20, B2 => lbl5_en1_n_133, Z => lbl5_en1_n_170);
  lbl5_en1_g6895 : AOI21D0BWP7T port map(A1 => lbl5_en1_n_155, A2 => FE_PHN225_lbl5_en1_new_period_4, B => lbl5_en1_n_142, ZN => lbl5_en1_n_169);
  lbl5_en1_g6896 : OAI211D1BWP7T port map(A1 => FE_PHN224_lbl5_en1_n_3, A2 => lbl5_en1_n_140, B => lbl5_en1_n_136, C => lbl5_en1_n_64, ZN => lbl5_en1_n_168);
  lbl5_en1_g6897 : AOI222D0BWP7T port map(A1 => lbl5_en1_n_141, A2 => FE_PHN221_lbl5_en1_new_period_14, B1 => lbl5_en1_n_115, B2 => lbl5_en1_n_98, C1 => lbl5_en1_n_58, C2 => direction_1(1), ZN => lbl5_en1_n_167);
  lbl5_en1_g6898 : MOAI22D0BWP7T port map(A1 => lbl5_en1_n_106, A2 => lbl5_en1_n_41, B1 => lbl5_en1_n_151, B2 => lbl5_en1_new_period(3), ZN => lbl5_en1_n_166);
  lbl5_en1_g6899 : IOA21D0BWP7T port map(A1 => lbl5_en1_n_140, A2 => lbl5_en1_n_126, B => FE_PHN216_lbl5_en1_new_period_8, ZN => lbl5_en1_n_164);
  lbl5_en1_g6900 : OAI31D0BWP7T port map(A1 => FE_PHN228_lbl5_en1_new_period_13, A2 => lbl5_en1_n_77, A3 => lbl5_en1_n_108, B => lbl5_en1_n_158, ZN => lbl5_en1_n_163);
  lbl5_en1_g6901 : OAI221D0BWP7T port map(A1 => lbl5_en1_n_106, A2 => lbl5_en1_n_22, B1 => lbl5_en1_n_21, B2 => lbl5_en1_n_108, C => lbl5_en1_n_154, ZN => lbl5_en1_n_165);
  lbl5_en1_g6903 : AOI21D0BWP7T port map(A1 => lbl5_en1_n_145, A2 => lbl5_en1_n_134, B => lbl5_en1_new_period(17), ZN => lbl5_en1_n_162);
  lbl5_en1_g6904 : OAI21D0BWP7T port map(A1 => lbl5_en1_n_108, A2 => FE_PHN203_lbl5_en1_new_period_15, B => lbl5_en1_n_154, ZN => lbl5_en1_n_161);
  lbl5_en1_g6905 : AO21D0BWP7T port map(A1 => lbl5_en1_n_58, A2 => direction_1(0), B => lbl5_en1_n_149, Z => lbl5_en1_n_160);
  lbl5_en1_g6907 : AOI221D0BWP7T port map(A1 => lbl5_en1_n_105, A2 => FE_PHN206_lbl5_en1_new_period_11, B1 => lbl5_en1_n_107, B2 => FE_PHN226_lbl5_en1_n_2, C => lbl5_en1_n_139, ZN => lbl5_en1_n_159);
  lbl5_en1_g6908 : OAI21D0BWP7T port map(A1 => lbl5_en1_n_128, A2 => lbl5_en1_n_103, B => FE_PHN228_lbl5_en1_new_period_13, ZN => lbl5_en1_n_158);
  lbl5_en1_g6909 : AO21D0BWP7T port map(A1 => lbl5_en1_n_109, A2 => FE_PHN321_lbl5_en1_new_period_1, B => lbl5_en1_n_144, Z => lbl5_en1_n_157);
  lbl5_en1_g6910 : AOI221D0BWP7T port map(A1 => lbl5_en1_n_105, A2 => FE_PHN250_lbl5_en1_new_period_5, B1 => lbl5_en1_n_107, B2 => FE_PHN245_lbl5_en1_n_10, C => lbl5_en1_n_147, ZN => lbl5_en1_n_156);
  lbl5_en1_g6911 : AO211D0BWP7T port map(A1 => lbl5_en1_n_107, A2 => lbl5_en1_n_41, B => lbl5_en1_n_144, C => lbl5_en1_n_110, Z => lbl5_en1_n_155);
  lbl5_en1_g6912 : INVD0BWP7T port map(I => lbl5_en1_n_154, ZN => lbl5_en1_n_153);
  lbl5_en1_g6913 : AOI221D0BWP7T port map(A1 => lbl5_en1_n_105, A2 => lbl5_en1_new_period(9), B1 => lbl5_en1_n_107, B2 => FE_PHN227_lbl5_en1_n_4, C => lbl5_en1_n_146, ZN => lbl5_en1_n_152);
  lbl5_en1_g6914 : AO21D0BWP7T port map(A1 => lbl5_en1_n_107, A2 => lbl5_en1_n_20, B => lbl5_en1_n_144, Z => lbl5_en1_n_151);
  lbl5_en1_g6915 : AO211D0BWP7T port map(A1 => lbl5_en1_n_111, A2 => FE_PHN211_lbl5_en1_new_period_0, B => lbl5_en1_n_118, C => lbl5_en0_rst, Z => lbl5_en1_n_150);
  lbl5_en1_g6916 : AOI21D0BWP7T port map(A1 => lbl5_en1_n_130, A2 => lbl5_en1_n_112, B => FE_PHN203_lbl5_en1_new_period_15, ZN => lbl5_en1_n_149);
  lbl5_en1_g6917 : AOI32D1BWP7T port map(A1 => lbl5_en1_n_120, A2 => lbl5_en1_n_7, A3 => FE_PHN206_lbl5_en1_new_period_11, B1 => lbl5_en1_n_105, B2 => lbl5_en1_n_78, ZN => lbl5_en1_n_148);
  lbl5_en1_g6918 : AOI211XD0BWP7T port map(A1 => lbl5_en1_n_105, A2 => FE_PHN221_lbl5_en1_new_period_14, B => lbl5_en1_n_141, C => lbl5_en1_n_115, ZN => lbl5_en1_n_154);
  lbl5_en1_g6919 : NR3D0BWP7T port map(A1 => lbl5_en1_n_117, A2 => lbl5_en1_n_20, A3 => lbl5_en1_new_period(3), ZN => lbl5_en1_n_143);
  lbl5_en1_g6920 : NR3D0BWP7T port map(A1 => lbl5_en1_n_117, A2 => lbl5_en1_n_41, A3 => FE_PHN225_lbl5_en1_new_period_4, ZN => lbl5_en1_n_142);
  lbl5_en1_g6921 : OAI221D0BWP7T port map(A1 => lbl5_en1_n_106, A2 => lbl5_en1_n_49, B1 => lbl5_en1_n_50, B2 => lbl5_en1_n_108, C => lbl5_en1_n_104, ZN => lbl5_en1_n_147);
  lbl5_en1_g6922 : OAI221D0BWP7T port map(A1 => lbl5_en1_n_106, A2 => lbl5_en1_n_67, B1 => lbl5_en1_n_66, B2 => lbl5_en1_n_108, C => lbl5_en1_n_104, ZN => lbl5_en1_n_146);
  lbl5_en1_g6923 : IND2D1BWP7T port map(A1 => lbl5_en1_n_130, B1 => lbl5_en1_n_22, ZN => lbl5_en1_n_145);
  lbl5_en1_g6924 : OAI221D0BWP7T port map(A1 => lbl5_en1_n_106, A2 => FE_PHN222_lbl5_en1_n_9, B1 => lbl5_crash_en, B2 => lbl5_en1_n_108, C => lbl5_en1_n_104, ZN => lbl5_en1_n_144);
  lbl5_en1_g6925 : ND3D0BWP7T port map(A1 => lbl5_en1_n_119, A2 => lbl5_en1_n_6, A3 => lbl5_en1_new_period(9), ZN => lbl5_en1_n_138);
  lbl5_en1_g6926 : IND3D1BWP7T port map(A1 => FE_PHN216_lbl5_en1_new_period_8, B1 => FE_PHN239_lbl5_en1_new_period_7, B2 => lbl5_en1_n_121, ZN => lbl5_en1_n_137);
  lbl5_en1_g6927 : IOA21D1BWP7T port map(A1 => lbl5_en1_n_116, A2 => lbl5_en1_n_122, B => FE_PHN224_lbl5_en1_n_3, ZN => lbl5_en1_n_136);
  lbl5_en1_g6928 : ND3D0BWP7T port map(A1 => lbl5_en1_n_123, A2 => FE_PHN223_lbl5_en1_n_8, A3 => FE_PHN250_lbl5_en1_new_period_5, ZN => lbl5_en1_n_135);
  lbl5_en1_g6929 : OAI221D0BWP7T port map(A1 => lbl5_en1_n_106, A2 => lbl5_en1_n_99, B1 => lbl5_en1_n_108, B2 => lbl5_en1_n_98, C => lbl5_en1_n_104, ZN => lbl5_en1_n_141);
  lbl5_en1_g6930 : AOI221D0BWP7T port map(A1 => lbl5_en1_n_105, A2 => lbl5_en1_n_57, B1 => lbl5_en1_n_107, B2 => lbl5_en1_n_56, C => lbl5_en1_n_103, ZN => lbl5_en1_n_140);
  lbl5_en1_g6931 : OAI221D0BWP7T port map(A1 => lbl5_en1_n_106, A2 => lbl5_en1_n_70, B1 => lbl5_en1_n_69, B2 => lbl5_en1_n_108, C => lbl5_en1_n_104, ZN => lbl5_en1_n_139);
  lbl5_en1_g6933 : IND2D1BWP7T port map(A1 => lbl5_en1_n_123, B1 => lbl5_en1_n_124, ZN => lbl5_en1_n_132);
  lbl5_en1_g6934 : IND2D1BWP7T port map(A1 => lbl5_en1_n_119, B1 => lbl5_en1_n_125, ZN => lbl5_en1_n_131);
  lbl5_en1_g6935 : IND2D1BWP7T port map(A1 => lbl5_en1_n_112, B1 => lbl5_en1_n_21, ZN => lbl5_en1_n_134);
  lbl5_en1_g6936 : IND2D1BWP7T port map(A1 => lbl5_en1_n_118, B1 => lbl5_en1_n_117, ZN => lbl5_en1_n_133);
  lbl5_en1_g6937 : NR2D0BWP7T port map(A1 => lbl5_en1_n_112, A2 => FE_PHN213_lbl5_en1_new_period_16, ZN => lbl5_en1_n_129);
  lbl5_en1_g6938 : MOAI22D0BWP7T port map(A1 => lbl5_en1_n_106, A2 => lbl5_en1_n_78, B1 => lbl5_en1_n_107, B2 => lbl5_en1_n_77, ZN => lbl5_en1_n_128);
  lbl5_en1_g6939 : IND2D1BWP7T port map(A1 => lbl5_en1_n_120, B1 => lbl5_en1_n_114, ZN => lbl5_en1_n_127);
  lbl5_en1_g6940 : AOI22D0BWP7T port map(A1 => lbl5_en1_n_105, A2 => FE_PHN239_lbl5_en1_new_period_7, B1 => lbl5_en1_n_107, B2 => lbl5_en1_n_3, ZN => lbl5_en1_n_126);
  lbl5_en1_g6941 : IND2D1BWP7T port map(A1 => FE_PHN221_lbl5_en1_new_period_14, B1 => lbl5_en1_n_113, ZN => lbl5_en1_n_130);
  lbl5_en1_g6942 : INVD1BWP7T port map(I => lbl5_en1_n_121, ZN => lbl5_en1_n_122);
  lbl5_en1_g6943 : ND2D1BWP7T port map(A1 => lbl5_en1_n_105, A2 => lbl5_en1_n_67, ZN => lbl5_en1_n_125);
  lbl5_en1_g6944 : ND2D1BWP7T port map(A1 => lbl5_en1_n_105, A2 => lbl5_en1_n_49, ZN => lbl5_en1_n_124);
  lbl5_en1_g6945 : INR2D1BWP7T port map(A1 => lbl5_en1_n_50, B1 => lbl5_en1_n_108, ZN => lbl5_en1_n_123);
  lbl5_en1_g6946 : NR2XD0BWP7T port map(A1 => lbl5_en1_n_108, A2 => lbl5_en1_n_56, ZN => lbl5_en1_n_121);
  lbl5_en1_g6947 : INR2D1BWP7T port map(A1 => lbl5_en1_n_69, B1 => lbl5_en1_n_108, ZN => lbl5_en1_n_120);
  lbl5_en1_g6948 : INR2D1BWP7T port map(A1 => lbl5_en1_n_66, B1 => lbl5_en1_n_108, ZN => lbl5_en1_n_119);
  lbl5_en1_g6949 : NR2D1BWP7T port map(A1 => lbl5_en1_n_106, A2 => FE_PHN211_lbl5_en1_new_period_0, ZN => lbl5_en1_n_118);
  lbl5_en1_g6950 : ND2D1BWP7T port map(A1 => lbl5_en1_n_107, A2 => lbl5_crash_en, ZN => lbl5_en1_n_117);
  lbl5_en1_g6951 : ND2D0BWP7T port map(A1 => lbl5_en1_n_108, A2 => lbl5_en1_n_104, ZN => lbl5_en1_n_111);
  lbl5_en1_g6952 : NR2D0BWP7T port map(A1 => lbl5_en1_n_106, A2 => lbl5_en1_n_42, ZN => lbl5_en1_n_110);
  lbl5_en1_g6953 : ND2D0BWP7T port map(A1 => lbl5_en1_n_106, A2 => lbl5_en1_n_108, ZN => lbl5_en1_n_109);
  lbl5_en1_g6954 : IND2D1BWP7T port map(A1 => lbl5_en1_n_57, B1 => lbl5_en1_n_105, ZN => lbl5_en1_n_116);
  lbl5_en1_g6955 : NR2D1BWP7T port map(A1 => lbl5_en1_n_108, A2 => FE_PHN221_lbl5_en1_new_period_14, ZN => lbl5_en1_n_115);
  lbl5_en1_g6956 : ND2D1BWP7T port map(A1 => lbl5_en1_n_105, A2 => lbl5_en1_n_70, ZN => lbl5_en1_n_114);
  lbl5_en1_g6957 : INR2D1BWP7T port map(A1 => lbl5_en1_n_99, B1 => lbl5_en1_n_106, ZN => lbl5_en1_n_113);
  lbl5_en1_g6958 : ND3D0BWP7T port map(A1 => lbl5_en1_n_107, A2 => lbl5_en1_n_98, A3 => FE_PHN221_lbl5_en1_new_period_14, ZN => lbl5_en1_n_112);
  lbl5_en1_g6959 : INVD1BWP7T port map(I => lbl5_en1_n_108, ZN => lbl5_en1_n_107);
  lbl5_en1_g6960 : IND4D0BWP7T port map(A1 => lbl5_engine_en, B1 => lbl5_en1_n_18, B2 => lbl5_en1_n_101, B3 => lbl5_en1_n_19, ZN => lbl5_en1_n_108);
  lbl5_en1_g6961 : INVD1BWP7T port map(I => lbl5_en1_n_106, ZN => lbl5_en1_n_105);
  lbl5_en1_g6962 : IND4D0BWP7T port map(A1 => lbl5_en1_n_60, B1 => lbl5_engine_en, B2 => lbl5_en1_n_18, B3 => lbl5_en1_n_101, ZN => lbl5_en1_n_106);
  lbl5_en1_g6963 : INVD0BWP7T port map(I => lbl5_en1_n_104, ZN => lbl5_en1_n_103);
  lbl5_en1_g6964 : ND2D1BWP7T port map(A1 => lbl5_en1_n_102, A2 => lbl5_en1_n_18, ZN => lbl5_en1_n_104);
  lbl5_en1_g6965 : NR2D1BWP7T port map(A1 => lbl5_en1_n_60, A2 => lbl5_en1_n_101, ZN => lbl5_en1_n_102);
  lbl5_en1_g6967 : NR4D0BWP7T port map(A1 => lbl5_en1_n_79, A2 => lbl5_en1_count(5), A3 => lbl5_en1_count(6), A4 => lbl5_en1_count(7), ZN => lbl5_en1_n_101);
  lbl5_en1_g6977 : AO221D0BWP7T port map(A1 => lbl5_en1_n_76, A2 => FE_PHN211_lbl5_en1_new_period_0, B1 => lbl5_en1_n_74, B2 => FE_PHN86_lbl5_en1_period_0, C => lbl5_en0_rst, Z => lbl5_en1_n_100);
  lbl5_en1_g7009 : MOAI22D0BWP7T port map(A1 => lbl5_en1_n_75, A2 => lbl5_en1_n_7, B1 => lbl5_en1_n_74, B2 => FE_PHN112_lbl5_en1_period_12, ZN => lbl5_en1_n_97);
  lbl5_en1_g7010 : AO22D0BWP7T port map(A1 => lbl5_en1_n_76, A2 => FE_PHN228_lbl5_en1_new_period_13, B1 => FE_PHN95_lbl5_en1_period_13, B2 => lbl5_en1_n_74, Z => lbl5_en1_n_96);
  lbl5_en1_g7011 : AO22D0BWP7T port map(A1 => lbl5_en1_n_76, A2 => lbl5_en1_new_period(18), B1 => FE_PHN87_lbl5_en1_period_18, B2 => lbl5_en1_n_74, Z => lbl5_en1_n_95);
  lbl5_en1_g7012 : MOAI22D0BWP7T port map(A1 => lbl5_en1_n_75, A2 => lbl5_en1_n_6, B1 => lbl5_en1_n_74, B2 => FE_PHN106_lbl5_en1_period_10, ZN => lbl5_en1_n_94);
  lbl5_en1_g7013 : AO22D0BWP7T port map(A1 => lbl5_en1_n_76, A2 => FE_PHN321_lbl5_en1_new_period_1, B1 => FE_PHN99_lbl5_en1_period_1, B2 => lbl5_en1_n_74, Z => lbl5_en1_n_93);
  lbl5_en1_g7014 : AO22D0BWP7T port map(A1 => lbl5_en1_n_76, A2 => FE_PHN244_lbl5_en1_new_period_2, B1 => FE_PHN70_lbl5_en1_period_2, B2 => lbl5_en1_n_74, Z => lbl5_en1_n_92);
  lbl5_en1_g7015 : AO22D0BWP7T port map(A1 => lbl5_en1_n_76, A2 => FE_PHN347_lbl5_en1_new_period_3, B1 => FE_PHN66_lbl5_en1_period_3, B2 => lbl5_en1_n_74, Z => lbl5_en1_n_91);
  lbl5_en1_g7016 : AO22D0BWP7T port map(A1 => lbl5_en1_n_76, A2 => FE_PHN225_lbl5_en1_new_period_4, B1 => FE_PHN147_lbl5_en1_period_4, B2 => lbl5_en1_n_74, Z => lbl5_en1_n_90);
  lbl5_en1_g7017 : MOAI22D0BWP7T port map(A1 => lbl5_en1_n_75, A2 => FE_PHN346_lbl5_en1_n_10, B1 => lbl5_en1_n_74, B2 => FE_PHN119_lbl5_en1_period_5, ZN => lbl5_en1_n_89);
  lbl5_en1_g7018 : MOAI22D0BWP7T port map(A1 => lbl5_en1_n_75, A2 => FE_PHN224_lbl5_en1_n_3, B1 => lbl5_en1_n_74, B2 => FE_PHN113_lbl5_en1_period_7, ZN => lbl5_en1_n_88);
  lbl5_en1_g7019 : MOAI22D0BWP7T port map(A1 => lbl5_en1_n_75, A2 => FE_PHN226_lbl5_en1_n_2, B1 => lbl5_en1_n_74, B2 => FE_PHN102_lbl5_en1_period_11, ZN => lbl5_en1_n_87);
  lbl5_en1_g7020 : MOAI22D0BWP7T port map(A1 => lbl5_en1_n_75, A2 => FE_PHN146_lbl5_en1_n_5, B1 => lbl5_en1_n_74, B2 => lbl5_en1_period(17), ZN => lbl5_en1_n_86);
  lbl5_en1_g7021 : AO22D0BWP7T port map(A1 => lbl5_en1_n_76, A2 => FE_PHN317_lbl5_en1_new_period_14, B1 => FE_PHN90_lbl5_en1_period_14, B2 => lbl5_en1_n_74, Z => lbl5_en1_n_85);
  lbl5_en1_g7022 : AO22D0BWP7T port map(A1 => lbl5_en1_n_76, A2 => FE_PHN203_lbl5_en1_new_period_15, B1 => FE_PHN84_lbl5_en1_period_15, B2 => lbl5_en1_n_74, Z => lbl5_en1_n_84);
  lbl5_en1_g7023 : MOAI22D0BWP7T port map(A1 => lbl5_en1_n_75, A2 => FE_PHN223_lbl5_en1_n_8, B1 => lbl5_en1_n_74, B2 => FE_PHN123_lbl5_en1_period_6, ZN => lbl5_en1_n_83);
  lbl5_en1_g7024 : AO22D0BWP7T port map(A1 => lbl5_en1_n_76, A2 => FE_PHN213_lbl5_en1_new_period_16, B1 => FE_PHN259_lbl5_en1_period_16, B2 => lbl5_en1_n_74, Z => lbl5_en1_n_82);
  lbl5_en1_g7025 : AO22D0BWP7T port map(A1 => lbl5_en1_n_76, A2 => FE_PHN312_lbl5_en1_new_period_8, B1 => FE_PHN89_lbl5_en1_period_8, B2 => lbl5_en1_n_74, Z => lbl5_en1_n_81);
  lbl5_en1_g7026 : MOAI22D0BWP7T port map(A1 => lbl5_en1_n_75, A2 => FE_PHN227_lbl5_en1_n_4, B1 => lbl5_en1_n_74, B2 => FE_PHN114_lbl5_en1_period_9, ZN => lbl5_en1_n_80);
  lbl5_en1_g7027 : INR2XD0BWP7T port map(A1 => lbl5_en1_n_78, B1 => FE_PHN228_lbl5_en1_new_period_13, ZN => lbl5_en1_n_99);
  lbl5_en1_g7028 : INR2XD0BWP7T port map(A1 => FE_PHN228_lbl5_en1_new_period_13, B1 => lbl5_en1_n_77, ZN => lbl5_en1_n_98);
  lbl5_en1_g7031 : IND3D1BWP7T port map(A1 => lbl5_en1_count(4), B1 => lbl5_en1_n_13, B2 => lbl5_en1_n_71, ZN => lbl5_en1_n_79);
  lbl5_en1_g7032 : AN3D1BWP7T port map(A1 => lbl5_en1_n_70, A2 => lbl5_en1_n_7, A3 => FE_PHN226_lbl5_en1_n_2, Z => lbl5_en1_n_78);
  lbl5_en1_g7033 : ND3D0BWP7T port map(A1 => lbl5_en1_n_69, A2 => lbl5_en1_new_period(12), A3 => FE_PHN206_lbl5_en1_new_period_11, ZN => lbl5_en1_n_77);
  lbl5_en1_g7034 : INVD1BWP7T port map(I => lbl5_en1_n_76, ZN => lbl5_en1_n_75);
  lbl5_en1_g7035 : NR2XD0BWP7T port map(A1 => lbl5_en0_rst, A2 => lbl5_en1_n_72, ZN => lbl5_en1_n_76);
  lbl5_en1_g7036 : NR2XD1BWP7T port map(A1 => lbl5_en0_rst, A2 => lbl5_en1_n_73, ZN => lbl5_en1_n_74);
  lbl5_en1_g7037 : INVD0BWP7T port map(I => lbl5_en1_n_73, ZN => lbl5_en1_n_72);
  lbl5_en1_g7038 : NR4D0BWP7T port map(A1 => lbl5_en1_n_61, A2 => lbl5_en1_count(3), A3 => lbl5_en1_count(2), A4 => lbl5_en1_count(1), ZN => lbl5_en1_n_71);
  lbl5_en1_g7039 : AOI211XD0BWP7T port map(A1 => lbl5_en1_n_319, A2 => lbl5_en1_n_14, B => lbl5_en1_n_68, C => lbl5_en1_n_17, ZN => lbl5_en1_n_73);
  lbl5_en1_g7040 : AN3D1BWP7T port map(A1 => lbl5_en1_n_67, A2 => lbl5_en1_n_6, A3 => FE_PHN227_lbl5_en1_n_4, Z => lbl5_en1_n_70);
  lbl5_en1_g7041 : AN3D1BWP7T port map(A1 => lbl5_en1_n_66, A2 => lbl5_en1_new_period(10), A3 => lbl5_en1_new_period(9), Z => lbl5_en1_n_69);
  lbl5_en1_g7042 : IND4D0BWP7T port map(A1 => lbl5_en1_n_54, B1 => lbl5_en1_n_29, B2 => lbl5_en1_n_45, B3 => lbl5_en1_n_62, ZN => lbl5_en1_n_68);
  lbl5_en1_g7043 : NR3D0BWP7T port map(A1 => lbl5_en1_n_57, A2 => FE_PHN239_lbl5_en1_new_period_7, A3 => FE_PHN216_lbl5_en1_new_period_8, ZN => lbl5_en1_n_67);
  lbl5_en1_g7044 : NR3D0BWP7T port map(A1 => lbl5_en1_n_56, A2 => lbl5_en1_n_11, A3 => FE_PHN224_lbl5_en1_n_3, ZN => lbl5_en1_n_66);
  lbl5_en1_g7045 : INVD1BWP7T port map(I => lbl5_en1_n_63, ZN => lbl5_en1_n_64);
  lbl5_en1_g7046 : NR2D1BWP7T port map(A1 => lbl5_en1_n_60, A2 => lbl5_en1_n_18, ZN => lbl5_en1_n_65);
  lbl5_en1_g7047 : IAO21D0BWP7T port map(A1 => lbl5_beep_en, A2 => lbl5_en1_n_55, B => lbl5_en0_rst, ZN => lbl5_en1_n_63);
  lbl5_en1_g7048 : NR4D0BWP7T port map(A1 => lbl5_en1_n_52, A2 => lbl5_en1_n_48, A3 => lbl5_en1_n_40, A4 => lbl5_en1_n_38, ZN => lbl5_en1_n_62);
  lbl5_en1_g7049 : OAI21D0BWP7T port map(A1 => lbl5_en1_n_53, A2 => lbl5_en1_frozen_boost, B => lbl5_en1_n_51, ZN => lbl5_en1_n_61);
  lbl5_en1_g7050 : INVD0BWP7T port map(I => lbl5_en1_n_59, ZN => lbl5_en1_n_58);
  lbl5_en1_g7051 : IND2D1BWP7T port map(A1 => lbl5_en1_n_55, B1 => lbl5_en1_n_19, ZN => lbl5_en1_n_60);
  lbl5_en1_g7052 : ND2D1BWP7T port map(A1 => lbl5_en1_n_19, A2 => lbl5_en1_n_55, ZN => lbl5_en1_n_59);
  lbl5_en1_g7053 : ND3D0BWP7T port map(A1 => lbl5_en1_n_49, A2 => FE_PHN223_lbl5_en1_n_8, A3 => FE_PHN245_lbl5_en1_n_10, ZN => lbl5_en1_n_57);
  lbl5_en1_g7054 : ND3D0BWP7T port map(A1 => lbl5_en1_n_50, A2 => lbl5_en1_new_period(6), A3 => FE_PHN250_lbl5_en1_new_period_5, ZN => lbl5_en1_n_56);
  lbl5_en1_g7055 : OAI211D1BWP7T port map(A1 => lbl5_en1_count(0), A2 => lbl5_en1_n_0, B => lbl5_en1_n_47, C => lbl5_en1_n_25, ZN => lbl5_en1_n_54);
  lbl5_en1_g7056 : AOI31D0BWP7T port map(A1 => lbl5_en1_n_26, A2 => lbl5_en1_n_24, A3 => lbl5_en1_prev_engine, B => lbl5_en1_n_16, ZN => lbl5_en1_n_55);
  lbl5_en1_g7057 : AOI21D0BWP7T port map(A1 => lbl5_en1_n_43, A2 => lbl5_en1_n_14, B => lbl5_en1_count(8), ZN => lbl5_en1_n_53);
  lbl5_en1_g7058 : OAI21D0BWP7T port map(A1 => lbl5_en1_n_319, A2 => lbl5_en1_n_14, B => lbl5_en1_n_46, ZN => lbl5_en1_n_52);
  lbl5_en1_g7059 : ND3D0BWP7T port map(A1 => lbl5_en1_n_44, A2 => lbl5_en1_n_14, A3 => lbl5_en1_frozen_boost, ZN => lbl5_en1_n_51);
  lbl5_en1_g7060 : OAI211D1BWP7T port map(A1 => lbl5_en1_n_15, A2 => lbl5_en1_n_320, B => lbl5_en1_n_23, C => lbl5_en1_n_31, ZN => lbl5_en1_n_48);
  lbl5_en1_g7061 : INR3D0BWP7T port map(A1 => lbl5_crash_en, B1 => lbl5_en1_n_12, B2 => lbl5_en1_n_41, ZN => lbl5_en1_n_50);
  lbl5_en1_g7062 : INR3D0BWP7T port map(A1 => lbl5_en1_n_42, B1 => FE_PHN211_lbl5_en1_new_period_0, B2 => FE_PHN225_lbl5_en1_new_period_4, ZN => lbl5_en1_n_49);
  lbl5_en1_g7063 : AOI211XD0BWP7T port map(A1 => lbl5_en1_n_0, A2 => lbl5_en1_count(0), B => lbl5_en1_n_35, C => lbl5_en1_n_30, ZN => lbl5_en1_n_47);
  lbl5_en1_g7064 : NR4D0BWP7T port map(A1 => lbl5_en1_n_34, A2 => lbl5_en1_n_39, A3 => lbl5_en1_n_36, A4 => lbl5_en1_n_28, ZN => lbl5_en1_n_46);
  lbl5_en1_g7065 : NR4D0BWP7T port map(A1 => lbl5_en1_n_33, A2 => lbl5_en1_n_37, A3 => lbl5_en1_n_32, A4 => lbl5_en1_n_27, ZN => lbl5_en1_n_45);
  lbl5_en1_g7066 : AOI31D0BWP7T port map(A1 => lbl5_en1_count(13), A2 => lbl5_en1_count(15), A3 => lbl5_en1_count(14), B => lbl5_en1_count(16), ZN => lbl5_en1_n_44);
  lbl5_en1_g7067 : AOI31D0BWP7T port map(A1 => lbl5_en1_count(15), A2 => lbl5_en1_count(16), A3 => lbl5_en1_count(14), B => lbl5_en1_count(18), ZN => lbl5_en1_n_43);
  lbl5_en1_g7068 : CKXOR2D1BWP7T port map(A1 => lbl5_en1_n_310, A2 => lbl5_en1_count(8), Z => lbl5_en1_n_40);
  lbl5_en1_g7069 : CKXOR2D1BWP7T port map(A1 => lbl5_en1_n_315, A2 => lbl5_en1_count(13), Z => lbl5_en1_n_39);
  lbl5_en1_g7070 : CKXOR2D1BWP7T port map(A1 => lbl5_en1_n_313, A2 => lbl5_en1_count(11), Z => lbl5_en1_n_38);
  lbl5_en1_g7071 : CKXOR2D1BWP7T port map(A1 => lbl5_en1_n_307, A2 => lbl5_en1_count(5), Z => lbl5_en1_n_37);
  lbl5_en1_g7072 : CKXOR2D1BWP7T port map(A1 => lbl5_en1_n_316, A2 => lbl5_en1_count(14), Z => lbl5_en1_n_36);
  lbl5_en1_g7073 : CKXOR2D1BWP7T port map(A1 => lbl5_en1_n_304, A2 => lbl5_en1_count(2), Z => lbl5_en1_n_35);
  lbl5_en1_g7074 : CKXOR2D1BWP7T port map(A1 => lbl5_en1_n_314, A2 => lbl5_en1_count(12), Z => lbl5_en1_n_34);
  lbl5_en1_g7076 : INR2XD0BWP7T port map(A1 => lbl5_en1_n_20, B1 => lbl5_en1_new_period(3), ZN => lbl5_en1_n_42);
  lbl5_en1_g7077 : IND2D1BWP7T port map(A1 => lbl5_en1_n_20, B1 => lbl5_en1_new_period(3), ZN => lbl5_en1_n_41);
  lbl5_en1_g7078 : CKXOR2D1BWP7T port map(A1 => lbl5_en1_n_306, A2 => lbl5_en1_count(4), Z => lbl5_en1_n_33);
  lbl5_en1_g7079 : CKXOR2D1BWP7T port map(A1 => lbl5_en1_n_309, A2 => lbl5_en1_count(7), Z => lbl5_en1_n_32);
  lbl5_en1_g7080 : XNR2D1BWP7T port map(A1 => lbl5_en1_n_312, A2 => lbl5_en1_count(10), ZN => lbl5_en1_n_31);
  lbl5_en1_g7081 : CKXOR2D1BWP7T port map(A1 => lbl5_en1_n_303, A2 => lbl5_en1_count(1), Z => lbl5_en1_n_30);
  lbl5_en1_g7082 : XNR2D1BWP7T port map(A1 => lbl5_en1_n_318, A2 => lbl5_en1_count(16), ZN => lbl5_en1_n_29);
  lbl5_en1_g7083 : CKXOR2D1BWP7T port map(A1 => lbl5_en1_n_317, A2 => lbl5_en1_count(15), Z => lbl5_en1_n_28);
  lbl5_en1_g7084 : CKXOR2D1BWP7T port map(A1 => lbl5_en1_n_308, A2 => lbl5_en1_count(6), Z => lbl5_en1_n_27);
  lbl5_en1_g7085 : MOAI22D0BWP7T port map(A1 => direction_1(1), A2 => lbl5_en1_prev_dir(1), B1 => direction_1(1), B2 => lbl5_en1_prev_dir(1), ZN => lbl5_en1_n_26);
  lbl5_en1_g7086 : XNR2D1BWP7T port map(A1 => lbl5_en1_n_305, A2 => lbl5_en1_count(3), ZN => lbl5_en1_n_25);
  lbl5_en1_g7087 : MOAI22D0BWP7T port map(A1 => direction_1(0), A2 => lbl5_en1_prev_dir(0), B1 => direction_1(0), B2 => lbl5_en1_prev_dir(0), ZN => lbl5_en1_n_24);
  lbl5_en1_g7088 : XNR2D1BWP7T port map(A1 => lbl5_en1_n_311, A2 => lbl5_en1_count(9), ZN => lbl5_en1_n_23);
  lbl5_en1_g7089 : NR2XD0BWP7T port map(A1 => FE_PHN213_lbl5_en1_new_period_16, A2 => FE_PHN203_lbl5_en1_new_period_15, ZN => lbl5_en1_n_22);
  lbl5_en1_g7090 : CKAN2D1BWP7T port map(A1 => FE_PHN213_lbl5_en1_new_period_16, A2 => FE_PHN203_lbl5_en1_new_period_15, Z => lbl5_en1_n_21);
  lbl5_en1_g7091 : NR2XD0BWP7T port map(A1 => FE_PHN348_lbl5_en1_new_period_1, A2 => FE_PHN244_lbl5_en1_new_period_2, ZN => lbl5_en1_n_20);
  lbl5_en1_g7092 : AN2D0BWP7T port map(A1 => lbl5_en1_n_320, A2 => lbl5_en1_n_15, Z => lbl5_en1_n_17);
  lbl5_en1_g7093 : NR2D1BWP7T port map(A1 => lbl5_en0_rst, A2 => lbl5_beep_en, ZN => lbl5_en1_n_19);
  lbl5_en1_g7094 : IND2D1BWP7T port map(A1 => lbl5_en1_prev_crash, B1 => lbl5_crash_en, ZN => lbl5_en1_n_18);
  lbl5_en1_g7095 : INVD0BWP7T port map(I => lbl5_engine_en, ZN => lbl5_en1_n_16);
  lbl5_en1_count_reg_0 : DFKCND1BWP7T port map(CN => FE_PHN117_lbl5_en1_n_13, CP => CTS_19, D => lbl5_en1_n_74, Q => lbl5_en1_count(0), QN => lbl5_en1_n_13);
  lbl5_en1_count_reg_17 : DFKCND1BWP7T port map(CN => lbl5_en1_n_74, CP => CTS_19, D => FE_PHN344_lbl5_en1_n_301, Q => lbl5_en1_count(17), QN => lbl5_en1_n_14);
  lbl5_en1_count_reg_18 : DFKCND1BWP7T port map(CN => lbl5_en1_n_74, CP => CTS_19, D => lbl5_en1_n_302, Q => lbl5_en1_count(18), QN => lbl5_en1_n_15);
  lbl5_en1_new_period_reg_0 : DFD1BWP7T port map(CP => CTS_20, D => lbl5_en1_n_150, Q => lbl5_en1_new_period(0), QN => lbl5_en1_n_9);
  lbl5_en1_new_period_reg_4 : DFD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_181, Q => lbl5_en1_new_period(4), QN => lbl5_en1_n_12);
  lbl5_en1_new_period_reg_5 : DFXD1BWP7T port map(CP => CTS_19, DA => lbl5_en1_n_147, DB => lbl5_en1_n_132, Q => lbl5_en1_new_period(5), QN => lbl5_en1_n_10, SA => FE_PHN345_lbl5_en1_new_period_5);
  lbl5_en1_new_period_reg_6 : DFD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_175, Q => lbl5_en1_new_period(6), QN => lbl5_en1_n_8);
  lbl5_en1_new_period_reg_7 : DFD1BWP7T port map(CP => CTS_20, D => lbl5_en1_n_168, Q => lbl5_en1_new_period(7), QN => lbl5_en1_n_3);
  lbl5_en1_new_period_reg_8 : DFD1BWP7T port map(CP => CTS_21, D => lbl5_en1_n_182, Q => lbl5_en1_new_period(8), QN => lbl5_en1_n_11);
  lbl5_en1_new_period_reg_9 : DFXD1BWP7T port map(CP => CTS_19, DA => lbl5_en1_n_146, DB => lbl5_en1_n_131, Q => FE_PHN215_lbl5_en1_new_period_9, QN => lbl5_en1_n_4, SA => lbl5_en1_new_period(9));
  lbl5_en1_new_period_reg_10 : DFD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_176, Q => lbl5_en1_new_period(10), QN => FE_PHN209_lbl5_en1_n_6);
  lbl5_en1_new_period_reg_11 : DFXD1BWP7T port map(CP => CTS_19, DA => lbl5_en1_n_139, DB => lbl5_en1_n_127, Q => lbl5_en1_new_period(11), QN => lbl5_en1_n_2, SA => FE_PHN206_lbl5_en1_new_period_11);
  lbl5_en1_new_period_reg_12 : DFD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_177, Q => lbl5_en1_new_period(12), QN => FE_PHN204_lbl5_en1_n_7);
  lbl5_en1_new_period_reg_17 : DFD1BWP7T port map(CP => CTS_19, D => lbl5_en1_n_180, Q => FE_PHN349_lbl5_en1_new_period_17, QN => lbl5_en1_n_5);
  lbl5_en1_g2 : MUX2ND0BWP7T port map(I0 => lbl5_en1_n_145, I1 => lbl5_en1_n_134, S => lbl5_en1_new_period(17), ZN => lbl5_en1_n_1);
  lbl5_en1_g7143 : MUX2ND0BWP7T port map(I0 => lbl5_en1_period(0), I1 => lbl5_en1_period(1), S => lbl5_en1_frozen_boost, ZN => lbl5_en1_n_0);
  lbl5_en1_g7144 : AO211D0BWP7T port map(A1 => lbl5_en1_n_276, A2 => lbl5_en1_n_275, B => lbl5_en1_n_202, C => lbl5_en1_n_277, Z => lbl5_en1_n_331);
  lbl5_en1_g7145 : OAI21D0BWP7T port map(A1 => lbl5_en1_n_236, A2 => lbl5_en1_n_264, B => lbl5_en1_n_216, ZN => lbl5_en1_n_332);
  lbl5_en1_frozen_boost_reg : DFXD1BWP7T port map(CP => CTS_19, DA => FE_PHN142_boost_audio_1, DB => FE_PHN140_lbl5_en1_frozen_boost, Q => lbl5_en1_frozen_boost, QN => lbl5_en1_n_282, SA => lbl5_en1_n_73);
  lbl5_en1_count_reg_16 : DFKCND1BWP7T port map(CN => lbl5_en1_n_74, CP => CTS_19, D => FE_PHN290_lbl5_en1_n_300, Q => lbl5_en1_count(16), QN => lbl5_en1_n_200);
  lbl5_en1_count_reg_13 : DFKCND1BWP7T port map(CN => lbl5_en1_n_74, CP => CTS_19, D => FE_PHN135_lbl5_en1_n_297, Q => lbl5_en1_count(13), QN => lbl5_en1_n_197);
  lbl5_en1_count_reg_15 : DFKCND1BWP7T port map(CN => lbl5_en1_n_74, CP => CTS_19, D => lbl5_en1_n_299, Q => lbl5_en1_count(15), QN => lbl5_en1_n_195);
  lbl5_en1_count_reg_12 : DFKCND1BWP7T port map(CN => FE_PHN148_lbl5_en1_n_296, CP => CTS_19, D => lbl5_en1_n_74, Q => lbl5_en1_count(12), QN => lbl5_en1_n_194);
  lbl5_en1_count_reg_7 : DFKCND1BWP7T port map(CN => FE_PHN159_lbl5_en1_n_291, CP => CTS_19, D => lbl5_en1_n_74, Q => lbl5_en1_count(7), QN => lbl5_en1_n_192);
  lbl5_en1_count_reg_11 : DFKCND1BWP7T port map(CN => lbl5_en1_n_295, CP => CTS_19, D => lbl5_en1_n_74, Q => lbl5_en1_count(11), QN => lbl5_en1_n_191);
  lbl5_en1_count_reg_14 : DFKCND1BWP7T port map(CN => lbl5_en1_n_74, CP => CTS_19, D => FE_PHN162_lbl5_en1_n_298, Q => lbl5_en1_count(14), QN => lbl5_en1_n_186);
  lbl5_en1_g7162 : IOA21D0BWP7T port map(A1 => lbl5_en1_n_319, A2 => lbl5_en1_n_195, B => lbl5_en1_count(14), ZN => lbl5_en1_n_333);
  lbl2_hscr_g18635 : IOA21D1BWP7T port map(A1 => lbl2_pixelator_color(3), A2 => lbl2_hscr_n_203, B => lbl2_hscr_n_370, ZN => lbl2_homescreen_color(3));
  lbl2_hscr_g18636 : IOA21D1BWP7T port map(A1 => lbl2_pixelator_color(2), A2 => lbl2_hscr_n_203, B => lbl2_hscr_n_370, ZN => lbl2_homescreen_color(2));
  lbl2_hscr_g18637 : IOA21D1BWP7T port map(A1 => lbl2_pixelator_color(1), A2 => lbl2_hscr_n_203, B => lbl2_hscr_n_371, ZN => lbl2_homescreen_color(1));
  lbl2_hscr_g18638 : IOA21D1BWP7T port map(A1 => lbl2_pixelator_color(0), A2 => lbl2_hscr_n_203, B => lbl2_hscr_n_371, ZN => lbl2_homescreen_color(0));
  lbl2_hscr_g18639 : IOA21D1BWP7T port map(A1 => lbl2_hscr_n_368, A2 => lbl2_hscr_n_345, B => lbl2_hscr_n_369, ZN => lbl2_hscr_n_371);
  lbl2_hscr_g18640 : IOA21D1BWP7T port map(A1 => lbl2_hscr_n_368, A2 => lbl2_hscr_n_328, B => lbl2_hscr_n_369, ZN => lbl2_hscr_n_370);
  lbl2_hscr_g18641 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_368, A2 => lbl2_hscr_n_360, B => lbl2_hscr_n_203, ZN => lbl2_hscr_n_369);
  lbl2_hscr_g18642 : AOI222D0BWP7T port map(A1 => lbl2_hscr_n_367, A2 => lbl2_hscr_n_180, B1 => lbl2_hscr_n_348, B2 => lbl2_hscr_n_32, C1 => lbl2_hscr_n_247, C2 => lbl2_hscr_n_110, ZN => lbl2_hscr_n_368);
  lbl2_hscr_g18643 : AOI211D1BWP7T port map(A1 => lbl2_hscr_n_10, A2 => lbl2_v_count(4), B => lbl2_hscr_n_366, C => lbl2_hscr_n_59, ZN => lbl2_hscr_n_367);
  lbl2_hscr_g18644 : OAI211D1BWP7T port map(A1 => lbl2_v_count(5), A2 => lbl2_hscr_n_10, B => lbl2_hscr_n_365, C => lbl2_hscr_n_38, ZN => lbl2_hscr_n_366);
  lbl2_hscr_g18645 : AO211D0BWP7T port map(A1 => lbl2_hscr_n_191, A2 => lbl2_hscr_n_198, B => lbl2_hscr_n_364, C => lbl2_hscr_n_291, Z => lbl2_hscr_n_365);
  lbl2_hscr_g18646 : IND4D0BWP7T port map(A1 => lbl2_hscr_n_363, B1 => lbl2_hscr_n_266, B2 => lbl2_hscr_n_344, B3 => lbl2_hscr_n_355, ZN => lbl2_hscr_n_364);
  lbl2_hscr_g18647 : ND4D0BWP7T port map(A1 => lbl2_hscr_n_362, A2 => lbl2_hscr_n_359, A3 => lbl2_hscr_n_361, A4 => lbl2_hscr_n_358, ZN => lbl2_hscr_n_363);
  lbl2_hscr_g18648 : OAI31D0BWP7T port map(A1 => lbl2_hscr_n_256, A2 => lbl2_hscr_n_321, A3 => lbl2_hscr_n_357, B => lbl2_h_count(0), ZN => lbl2_hscr_n_362);
  lbl2_hscr_g18649 : OAI31D0BWP7T port map(A1 => lbl2_hscr_n_210, A2 => lbl2_hscr_n_299, A3 => lbl2_hscr_n_350, B => FE_DBTN19_lbl2_h_count_1, ZN => lbl2_hscr_n_361);
  lbl2_hscr_g18650 : ND4D0BWP7T port map(A1 => lbl2_hscr_n_349, A2 => lbl2_hscr_n_73, A3 => lbl2_hscr_n_35, A4 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_360);
  lbl2_hscr_g18651 : NR4D0BWP7T port map(A1 => lbl2_hscr_n_352, A2 => lbl2_hscr_n_356, A3 => lbl2_hscr_n_343, A4 => lbl2_hscr_n_325, ZN => lbl2_hscr_n_359);
  lbl2_hscr_g18652 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_306, A2 => lbl2_hscr_n_103, B1 => lbl2_hscr_n_239, B2 => lbl2_hscr_n_71, C => lbl2_hscr_n_354, ZN => lbl2_hscr_n_358);
  lbl2_hscr_g18653 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_143, A2 => lbl2_hscr_n_209, B => lbl2_hscr_n_353, C => lbl2_hscr_n_212, ZN => lbl2_hscr_n_357);
  lbl2_hscr_g18654 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_351, A2 => FE_DBTN19_lbl2_h_count_1, ZN => lbl2_hscr_n_356);
  lbl2_hscr_g18655 : OAI31D0BWP7T port map(A1 => lbl2_hscr_n_257, A2 => lbl2_hscr_n_290, A3 => lbl2_hscr_n_341, B => lbl2_h_count(2), ZN => lbl2_hscr_n_355);
  lbl2_hscr_g18656 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_347, A2 => lbl2_h_count(2), B1 => lbl2_hscr_n_208, B2 => lbl2_hscr_n_138, ZN => lbl2_hscr_n_354);
  lbl2_hscr_g18657 : MAOI22D0BWP7T port map(A1 => lbl2_hscr_n_288, A2 => lbl2_hscr_n_103, B1 => lbl2_hscr_n_346, B2 => FE_DBTN19_lbl2_h_count_1, ZN => lbl2_hscr_n_353);
  lbl2_hscr_g18658 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_333, A2 => lbl2_hscr_n_300, A3 => lbl2_hscr_n_223, B => lbl2_h_count(0), ZN => lbl2_hscr_n_352);
  lbl2_hscr_g18659 : NR4D0BWP7T port map(A1 => lbl2_hscr_n_336, A2 => lbl2_hscr_n_321, A3 => lbl2_hscr_n_282, A4 => lbl2_hscr_n_256, ZN => lbl2_hscr_n_351);
  lbl2_hscr_g18660 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_82, A2 => lbl2_hscr_n_242, B => lbl2_hscr_n_342, C => lbl2_hscr_n_223, ZN => lbl2_hscr_n_350);
  lbl2_hscr_g18661 : MAOI22D0BWP7T port map(A1 => lbl2_hscr_n_51, A2 => lbl2_v_count(6), B1 => lbl2_hscr_n_345, B2 => lbl2_hscr_n_328, ZN => lbl2_hscr_n_349);
  lbl2_hscr_g18662 : AOI211D1BWP7T port map(A1 => lbl2_hscr_n_308, A2 => lbl2_hscr_n_6, B => lbl2_hscr_n_338, C => lbl2_hscr_n_58, ZN => lbl2_hscr_n_348);
  lbl2_hscr_g18663 : NR4D0BWP7T port map(A1 => lbl2_hscr_n_330, A2 => lbl2_hscr_n_302, A3 => lbl2_hscr_n_292, A4 => lbl2_hscr_n_270, ZN => lbl2_hscr_n_347);
  lbl2_hscr_g18664 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_273, A2 => FE_DBTN20_lbl2_h_count_2, B1 => lbl2_hscr_n_293, B2 => lbl2_hscr_n_156, C => lbl2_hscr_n_339, ZN => lbl2_hscr_n_346);
  lbl2_hscr_g18665 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_269, A2 => lbl2_hscr_n_116, B1 => lbl2_hscr_n_253, B2 => lbl2_v_count(1), C => lbl2_hscr_n_334, ZN => lbl2_hscr_n_344);
  lbl2_hscr_g18666 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_161, A2 => lbl2_hscr_n_244, B => lbl2_hscr_n_335, C => lbl2_hscr_n_276, ZN => lbl2_hscr_n_345);
  lbl2_hscr_g18667 : OA31D1BWP7T port map(A1 => lbl2_hscr_n_257, A2 => lbl2_hscr_n_283, A3 => lbl2_hscr_n_326, B => lbl2_hscr_n_29, Z => lbl2_hscr_n_343);
  lbl2_hscr_g18668 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_250, A2 => lbl2_hscr_n_120, B1 => lbl2_hscr_n_232, B2 => lbl2_hscr_n_133, C => lbl2_hscr_n_340, ZN => lbl2_hscr_n_342);
  lbl2_hscr_g18669 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_206, A2 => lbl2_hscr_n_47, B => lbl2_hscr_n_337, ZN => lbl2_hscr_n_341);
  lbl2_hscr_g18670 : OAI211D1BWP7T port map(A1 => lbl2_v_count(0), A2 => lbl2_hscr_n_233, B => lbl2_hscr_n_327, C => lbl2_hscr_n_296, ZN => lbl2_hscr_n_340);
  lbl2_hscr_g18671 : ND4D0BWP7T port map(A1 => lbl2_hscr_n_322, A2 => lbl2_hscr_n_286, A3 => lbl2_hscr_n_261, A4 => lbl2_hscr_n_260, ZN => lbl2_hscr_n_339);
  lbl2_hscr_g18672 : IND4D0BWP7T port map(A1 => lbl2_v_count(5), B1 => lbl2_v_count(8), B2 => lbl2_hscr_n_26, B3 => lbl2_hscr_n_320, ZN => lbl2_hscr_n_338);
  lbl2_hscr_g18673 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_317, A2 => lbl2_hscr_n_47, B1 => lbl2_hscr_n_168, B2 => lbl2_hscr_n_183, C => lbl2_hscr_n_210, ZN => lbl2_hscr_n_337);
  lbl2_hscr_g18674 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_123, A2 => lbl2_hscr_n_274, B => lbl2_hscr_n_323, C => lbl2_hscr_n_304, ZN => lbl2_hscr_n_336);
  lbl2_hscr_g18675 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_204, A2 => lbl2_hscr_n_198, A3 => lbl2_hscr_n_25, B => lbl2_hscr_n_331, ZN => lbl2_hscr_n_335);
  lbl2_hscr_g18676 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_226, A2 => lbl2_hscr_n_147, B => lbl2_hscr_n_329, C => lbl2_hscr_n_215, ZN => lbl2_hscr_n_334);
  lbl2_hscr_g18677 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_210, A2 => lbl2_v_count(0), B => lbl2_hscr_n_332, ZN => lbl2_hscr_n_333);
  lbl2_hscr_g18678 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_164, A2 => lbl2_hscr_n_200, B => lbl2_hscr_n_324, C => lbl2_hscr_n_211, ZN => lbl2_hscr_n_332);
  lbl2_hscr_g18679 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_315, A2 => lbl2_hscr_n_48, B => lbl2_hscr_n_316, ZN => lbl2_hscr_n_331);
  lbl2_hscr_g18680 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_298, A2 => lbl2_hscr_n_259, A3 => lbl2_hscr_n_255, B => lbl2_hscr_n_47, ZN => lbl2_hscr_n_330);
  lbl2_hscr_g18681 : AOI211XD0BWP7T port map(A1 => lbl2_hscr_n_163, A2 => lbl2_hscr_n_182, B => lbl2_hscr_n_313, C => lbl2_hscr_n_301, ZN => lbl2_hscr_n_329);
  lbl2_hscr_g18682 : OA221D0BWP7T port map(A1 => lbl2_hscr_n_207, A2 => lbl2_hscr_n_158, B1 => lbl2_hscr_n_142, B2 => lbl2_hscr_n_208, C => lbl2_hscr_n_314, Z => lbl2_hscr_n_327);
  lbl2_hscr_g18683 : OAI31D0BWP7T port map(A1 => lbl2_hscr_n_68, A2 => lbl2_hscr_n_145, A3 => lbl2_hscr_n_243, B => lbl2_hscr_n_319, ZN => lbl2_hscr_n_326);
  lbl2_hscr_g18684 : OAI221D0BWP7T port map(A1 => lbl2_hscr_n_271, A2 => lbl2_hscr_n_145, B1 => lbl2_hscr_n_91, B2 => lbl2_hscr_n_246, C => lbl2_hscr_n_318, ZN => lbl2_hscr_n_328);
  lbl2_hscr_g18685 : AOI211D1BWP7T port map(A1 => lbl2_hscr_n_305, A2 => lbl2_hscr_n_233, B => lbl2_h_count(1), C => lbl2_hscr_n_9, ZN => lbl2_hscr_n_325);
  lbl2_hscr_g18686 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_234, A2 => lbl2_hscr_n_103, A3 => lbl2_hscr_n_47, B1 => lbl2_hscr_n_309, B2 => lbl2_h_count(1), ZN => lbl2_hscr_n_324);
  lbl2_hscr_g18687 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_175, A2 => lbl2_hscr_n_116, A3 => lbl2_hscr_n_71, B1 => lbl2_hscr_n_310, B2 => lbl2_hscr_n_103, ZN => lbl2_hscr_n_323);
  lbl2_hscr_g18688 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_303, A2 => lbl2_h_count(2), B1 => lbl2_hscr_n_251, B2 => lbl2_hscr_n_122, ZN => lbl2_hscr_n_322);
  lbl2_hscr_g18689 : AOI211D1BWP7T port map(A1 => lbl2_v_count(2), A2 => lbl2_v_count(4), B => lbl2_hscr_n_311, C => lbl2_hscr_n_238, ZN => lbl2_hscr_n_320);
  lbl2_hscr_g18690 : OA221D0BWP7T port map(A1 => lbl2_hscr_n_200, A2 => lbl2_hscr_n_141, B1 => lbl2_hscr_n_121, B2 => lbl2_hscr_n_208, C => lbl2_hscr_n_307, Z => lbl2_hscr_n_319);
  lbl2_hscr_g18691 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_236, A2 => lbl2_hscr_n_192, B1 => lbl2_hscr_n_267, B2 => lbl2_hscr_n_159, C => lbl2_hscr_n_294, ZN => lbl2_hscr_n_318);
  lbl2_hscr_g18692 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_155, A2 => lbl2_hscr_n_184, B => lbl2_hscr_n_280, C => lbl2_hscr_n_264, ZN => lbl2_hscr_n_321);
  lbl2_hscr_g18693 : AO221D0BWP7T port map(A1 => lbl2_hscr_n_195, A2 => lbl2_hscr_n_159, B1 => lbl2_hscr_n_269, B2 => lbl2_hscr_n_64, C => lbl2_hscr_n_187, Z => lbl2_hscr_n_317);
  lbl2_hscr_g18694 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_275, A2 => lbl2_hscr_n_159, A3 => lbl2_hscr_n_48, B1 => lbl2_hscr_n_284, B2 => lbl2_hscr_n_180, ZN => lbl2_hscr_n_316);
  lbl2_hscr_g18695 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_221, A2 => lbl2_hscr_n_114, A3 => lbl2_hscr_n_116, B => lbl2_hscr_n_312, ZN => lbl2_hscr_n_315);
  lbl2_hscr_g18696 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_289, A2 => lbl2_hscr_n_71, B1 => lbl2_hscr_n_199, B2 => lbl2_hscr_n_169, ZN => lbl2_hscr_n_314);
  lbl2_hscr_g18697 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_295, A2 => lbl2_hscr_n_90, B1 => lbl2_hscr_n_262, B2 => lbl2_hscr_n_47, ZN => lbl2_hscr_n_313);
  lbl2_hscr_g18698 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_244, A2 => lbl2_hscr_n_64, B => lbl2_hscr_n_285, ZN => lbl2_hscr_n_312);
  lbl2_hscr_g18699 : OAI31D0BWP7T port map(A1 => direction_between(3), A2 => lbl2_hscr_n_66, A3 => lbl2_hscr_n_278, B => lbl2_hscr_n_150, ZN => lbl2_hscr_n_311);
  lbl2_hscr_g18700 : AO211D0BWP7T port map(A1 => lbl2_hscr_n_227, A2 => lbl2_hscr_n_98, B => lbl2_hscr_n_288, C => lbl2_hscr_n_224, Z => lbl2_hscr_n_310);
  lbl2_hscr_g18701 : OAI221D0BWP7T port map(A1 => lbl2_hscr_n_233, A2 => lbl2_hscr_n_2, B1 => lbl2_hscr_n_47, B2 => lbl2_hscr_n_255, C => lbl2_hscr_n_287, ZN => lbl2_hscr_n_309);
  lbl2_hscr_g18702 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_278, A2 => direction_between(2), B => lbl2_central_x_vec(8), ZN => lbl2_hscr_n_308);
  lbl2_hscr_g18703 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_194, A2 => lbl2_hscr_n_118, A3 => lbl2_hscr_n_71, B => lbl2_hscr_n_281, ZN => lbl2_hscr_n_307);
  lbl2_hscr_g18704 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_117, A2 => lbl2_hscr_n_229, B => lbl2_hscr_n_245, C => lbl2_hscr_n_265, ZN => lbl2_hscr_n_306);
  lbl2_hscr_g18705 : AOI222D0BWP7T port map(A1 => lbl2_hscr_n_199, A2 => lbl2_hscr_n_140, B1 => lbl2_hscr_n_250, B2 => lbl2_hscr_n_97, C1 => lbl2_hscr_n_254, C2 => lbl2_hscr_n_64, ZN => lbl2_hscr_n_305);
  lbl2_hscr_g18706 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_263, A2 => FE_DBTN20_lbl2_h_count_2, B1 => lbl2_hscr_n_199, B2 => lbl2_hscr_n_178, ZN => lbl2_hscr_n_304);
  lbl2_hscr_g18707 : AO21D0BWP7T port map(A1 => lbl2_hscr_n_182, A2 => lbl2_hscr_n_137, B => lbl2_hscr_n_297, Z => lbl2_hscr_n_303);
  lbl2_hscr_g18708 : OAI32D1BWP7T port map(A1 => lbl2_hscr_n_101, A2 => lbl2_hscr_n_134, A3 => lbl2_hscr_n_193, B1 => lbl2_hscr_n_96, B2 => lbl2_hscr_n_279, ZN => lbl2_hscr_n_302);
  lbl2_hscr_g18709 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_279, A2 => lbl2_hscr_n_124, B1 => lbl2_hscr_n_214, B2 => lbl2_v_count(1), ZN => lbl2_hscr_n_301);
  lbl2_hscr_g18710 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_277, A2 => lbl2_hscr_n_47, B1 => lbl2_hscr_n_250, B2 => lbl2_hscr_n_176, ZN => lbl2_hscr_n_300);
  lbl2_hscr_g18711 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_268, A2 => lbl2_hscr_n_91, B1 => lbl2_hscr_n_220, B2 => lbl2_hscr_n_48, ZN => lbl2_hscr_n_299);
  lbl2_hscr_g18712 : OA22D0BWP7T port map(A1 => lbl2_hscr_n_272, A2 => lbl2_hscr_n_161, B1 => lbl2_hscr_n_138, B2 => lbl2_hscr_n_226, Z => lbl2_hscr_n_298);
  lbl2_hscr_g18713 : AOI211D1BWP7T port map(A1 => lbl2_hscr_n_228, A2 => lbl2_hscr_n_229, B => lbl2_hscr_n_117, C => lbl2_hscr_n_82, ZN => lbl2_hscr_n_297);
  lbl2_hscr_g18714 : IND4D0BWP7T port map(A1 => lbl2_hscr_n_124, B1 => lbl2_h_count(2), B2 => lbl2_v_count(1), B3 => lbl2_hscr_n_227, ZN => lbl2_hscr_n_296);
  lbl2_hscr_g18715 : OA211D0BWP7T port map(A1 => lbl2_hscr_n_99, A2 => lbl2_hscr_n_226, B => lbl2_hscr_n_245, C => lbl2_hscr_n_222, Z => lbl2_hscr_n_295);
  lbl2_hscr_g18716 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_246, A2 => lbl2_hscr_n_116, A3 => lbl2_hscr_n_82, ZN => lbl2_hscr_n_294);
  lbl2_hscr_g18717 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_243, A2 => lbl2_hscr_n_83, B => lbl2_hscr_n_173, ZN => lbl2_hscr_n_293);
  lbl2_hscr_g18718 : AOI211D1BWP7T port map(A1 => lbl2_hscr_n_243, A2 => lbl2_hscr_n_173, B => lbl2_hscr_n_101, C => lbl2_hscr_n_145, ZN => lbl2_hscr_n_292);
  lbl2_hscr_g18719 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_242, A2 => lbl2_hscr_n_235, B => lbl2_hscr_n_91, ZN => lbl2_hscr_n_291);
  lbl2_hscr_g18720 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_242, A2 => lbl2_hscr_n_82, A3 => lbl2_hscr_n_83, ZN => lbl2_hscr_n_290);
  lbl2_hscr_g18721 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_234, B1 => lbl2_hscr_n_258, ZN => lbl2_hscr_n_289);
  lbl2_hscr_g18722 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_250, A2 => lbl2_hscr_n_140, B1 => lbl2_hscr_n_199, B2 => lbl2_hscr_n_97, ZN => lbl2_hscr_n_287);
  lbl2_hscr_g18723 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_225, A2 => lbl2_hscr_n_153, A3 => lbl2_hscr_n_67, B1 => lbl2_hscr_n_232, B2 => lbl2_hscr_n_144, ZN => lbl2_hscr_n_286);
  lbl2_hscr_g18724 : AOI33D1BWP7T port map(A1 => lbl2_hscr_n_204, A2 => lbl2_hscr_n_216, A3 => lbl2_hscr_n_145, B1 => lbl2_hscr_n_194, B2 => lbl2_hscr_n_180, B3 => lbl2_hscr_n_51, ZN => lbl2_hscr_n_285);
  lbl2_hscr_g18725 : OAI33D1BWP7T port map(A1 => lbl2_hscr_n_47, A2 => lbl2_hscr_n_116, A3 => lbl2_hscr_n_218, B1 => lbl2_hscr_n_52, B2 => lbl2_hscr_n_171, B3 => lbl2_hscr_n_155, ZN => lbl2_hscr_n_284);
  lbl2_hscr_g18726 : OAI33D1BWP7T port map(A1 => lbl2_hscr_n_1, A2 => lbl2_hscr_n_82, A3 => lbl2_hscr_n_213, B1 => FE_DBTN20_lbl2_h_count_2, B2 => lbl2_hscr_n_119, B3 => lbl2_hscr_n_229, ZN => lbl2_hscr_n_283);
  lbl2_hscr_g18727 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_209, A2 => lbl2_hscr_n_127, B1 => lbl2_hscr_n_249, B2 => lbl2_hscr_n_158, ZN => lbl2_hscr_n_282);
  lbl2_hscr_g18728 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_240, A2 => lbl2_hscr_n_230, B1 => lbl2_hscr_n_207, B2 => lbl2_hscr_n_148, ZN => lbl2_hscr_n_281);
  lbl2_hscr_g18729 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_250, A2 => lbl2_hscr_n_167, B1 => lbl2_hscr_n_232, B2 => lbl2_hscr_n_157, ZN => lbl2_hscr_n_280);
  lbl2_hscr_g18730 : OAI31D0BWP7T port map(A1 => lbl2_hscr_n_116, A2 => lbl2_hscr_n_135, A3 => lbl2_hscr_n_231, B => lbl2_hscr_n_235, ZN => lbl2_hscr_n_288);
  lbl2_hscr_g18731 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_230, A2 => lbl2_hscr_n_149, B => lbl2_hscr_n_220, ZN => lbl2_hscr_n_277);
  lbl2_hscr_g18732 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_230, B1 => lbl2_hscr_n_50, B2 => lbl2_hscr_n_180, ZN => lbl2_hscr_n_276);
  lbl2_hscr_g18733 : IOA21D1BWP7T port map(A1 => lbl2_hscr_n_221, A2 => lbl2_hscr_n_108, B => lbl2_hscr_n_217, ZN => lbl2_hscr_n_275);
  lbl2_hscr_g18734 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_183, A2 => lbl2_hscr_n_2, A3 => lbl2_h_count(2), B => lbl2_hscr_n_251, ZN => lbl2_hscr_n_274);
  lbl2_hscr_g18735 : OAI31D0BWP7T port map(A1 => lbl2_v_count(0), A2 => lbl2_hscr_n_101, A3 => lbl2_hscr_n_197, B => lbl2_hscr_n_252, ZN => lbl2_hscr_n_273);
  lbl2_hscr_g18736 : OA21D0BWP7T port map(A1 => lbl2_hscr_n_231, A2 => lbl2_hscr_n_104, B => lbl2_hscr_n_184, Z => lbl2_hscr_n_272);
  lbl2_hscr_g18737 : IND4D0BWP7T port map(A1 => lbl2_hscr_n_90, B1 => lbl2_hscr_n_76, B2 => lbl2_hscr_n_172, B3 => lbl2_hscr_n_205, ZN => lbl2_hscr_n_271);
  lbl2_hscr_g18738 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_228, A2 => lbl2_hscr_n_117, A3 => lbl2_hscr_n_1, ZN => lbl2_hscr_n_270);
  lbl2_hscr_g18739 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_226, A2 => lbl2_hscr_n_1, B => lbl2_hscr_n_202, ZN => lbl2_hscr_n_279);
  lbl2_hscr_g18740 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_9, A2 => lbl2_hscr_n_84, B => lbl2_hscr_n_248, C => lbl2_hscr_n_81, ZN => lbl2_hscr_n_278);
  lbl2_hscr_g18741 : INVD0BWP7T port map(I => lbl2_hscr_n_269, ZN => lbl2_hscr_n_268);
  lbl2_hscr_g18742 : AO22D0BWP7T port map(A1 => lbl2_hscr_n_236, A2 => lbl2_hscr_n_50, B1 => lbl2_hscr_n_108, B2 => lbl2_hscr_n_205, Z => lbl2_hscr_n_267);
  lbl2_hscr_g18743 : IOA21D1BWP7T port map(A1 => lbl2_hscr_n_138, A2 => lbl2_hscr_n_96, B => lbl2_hscr_n_251, ZN => lbl2_hscr_n_266);
  lbl2_hscr_g18744 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_231, A2 => lbl2_hscr_n_143, B => lbl2_hscr_n_241, ZN => lbl2_hscr_n_265);
  lbl2_hscr_g18745 : OA33D0BWP7T port map(A1 => lbl2_hscr_n_101, A2 => lbl2_hscr_n_172, A3 => lbl2_hscr_n_173, B1 => lbl2_v_count(1), B2 => lbl2_hscr_n_96, B3 => lbl2_hscr_n_201, Z => lbl2_hscr_n_264);
  lbl2_hscr_g18746 : OAI32D1BWP7T port map(A1 => lbl2_hscr_n_47, A2 => lbl2_hscr_n_134, A3 => lbl2_hscr_n_181, B1 => lbl2_hscr_n_124, B2 => lbl2_hscr_n_226, ZN => lbl2_hscr_n_263);
  lbl2_hscr_g18747 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_202, A2 => lbl2_hscr_n_137, B => lbl2_hscr_n_253, ZN => lbl2_hscr_n_262);
  lbl2_hscr_g18748 : OA22D0BWP7T port map(A1 => lbl2_hscr_n_237, A2 => lbl2_hscr_n_90, B1 => lbl2_hscr_n_48, B2 => lbl2_hscr_n_206, Z => lbl2_hscr_n_261);
  lbl2_hscr_g18749 : OA22D0BWP7T port map(A1 => lbl2_hscr_n_222, A2 => lbl2_hscr_n_102, B1 => lbl2_hscr_n_96, B2 => lbl2_hscr_n_209, Z => lbl2_hscr_n_260);
  lbl2_hscr_g18750 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_0, A2 => lbl2_hscr_n_82, B1 => lbl2_hscr_n_202, B2 => lbl2_hscr_n_122, ZN => lbl2_hscr_n_259);
  lbl2_hscr_g18751 : MAOI22D0BWP7T port map(A1 => lbl2_hscr_n_227, A2 => lbl2_hscr_n_118, B1 => lbl2_hscr_n_154, B2 => lbl2_hscr_n_142, ZN => lbl2_hscr_n_258);
  lbl2_hscr_g18752 : OAI22D0BWP7T port map(A1 => lbl2_hscr_n_193, A2 => lbl2_hscr_n_125, B1 => lbl2_hscr_n_229, B2 => lbl2_hscr_n_106, ZN => lbl2_hscr_n_269);
  lbl2_hscr_g18753 : INVD0BWP7T port map(I => lbl2_hscr_n_255, ZN => lbl2_hscr_n_254);
  lbl2_hscr_g18754 : INVD0BWP7T port map(I => lbl2_hscr_n_252, ZN => lbl2_hscr_n_253);
  lbl2_hscr_g18755 : INVD0BWP7T port map(I => lbl2_hscr_n_250, ZN => lbl2_hscr_n_249);
  lbl2_hscr_g18756 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_126, A2 => lbl2_h_count(2), B => lbl2_hscr_n_219, ZN => lbl2_hscr_n_248);
  lbl2_hscr_g18757 : OAI31D0BWP7T port map(A1 => lbl2_h_count(4), A2 => lbl2_h_count(2), A3 => lbl2_hscr_n_177, B => lbl2_hscr_n_185, ZN => lbl2_hscr_n_247);
  lbl2_hscr_g18758 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_170, A2 => lbl2_hscr_n_228, ZN => lbl2_hscr_n_257);
  lbl2_hscr_g18759 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_190, A2 => lbl2_hscr_n_47, A3 => lbl2_h_count(2), ZN => lbl2_hscr_n_256);
  lbl2_hscr_g18760 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_231, B1 => lbl2_hscr_n_137, ZN => lbl2_hscr_n_255);
  lbl2_hscr_g18761 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_226, B1 => lbl2_hscr_n_118, ZN => lbl2_hscr_n_252);
  lbl2_hscr_g18762 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_226, A2 => lbl2_hscr_n_64, ZN => lbl2_hscr_n_251);
  lbl2_hscr_g18763 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_230, A2 => FE_DBTN20_lbl2_h_count_2, ZN => lbl2_hscr_n_250);
  lbl2_hscr_g18764 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_123, A2 => lbl2_hscr_n_121, B => lbl2_hscr_n_226, ZN => lbl2_hscr_n_241);
  lbl2_hscr_g18765 : OA221D0BWP7T port map(A1 => lbl2_hscr_n_117, A2 => lbl2_hscr_n_12, B1 => lbl2_hscr_n_1, B2 => lbl2_hscr_n_141, C => lbl2_hscr_n_188, Z => lbl2_hscr_n_240);
  lbl2_hscr_g18766 : OAI31D0BWP7T port map(A1 => lbl2_hscr_n_64, A2 => lbl2_hscr_n_172, A3 => lbl2_hscr_n_174, B => lbl2_hscr_n_206, ZN => lbl2_hscr_n_239);
  lbl2_hscr_g18767 : OAI211D1BWP7T port map(A1 => lbl2_v_count(2), A2 => lbl2_hscr_n_30, B => lbl2_hscr_n_189, C => lbl2_hscr_n_151, ZN => lbl2_hscr_n_238);
  lbl2_hscr_g18768 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_55, A2 => lbl2_hscr_n_54, B => lbl2_hscr_n_205, C => lbl2_hscr_n_172, ZN => lbl2_hscr_n_246);
  lbl2_hscr_g18769 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_160, A2 => lbl2_hscr_n_133, A3 => lbl2_hscr_n_145, B1 => lbl2_hscr_n_202, B2 => lbl2_hscr_n_98, ZN => lbl2_hscr_n_245);
  lbl2_hscr_g18770 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_204, A2 => lbl2_hscr_n_172, A3 => lbl2_hscr_n_50, ZN => lbl2_hscr_n_244);
  lbl2_hscr_g18771 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_195, A2 => lbl2_v_count(1), A3 => lbl2_v_count(0), ZN => lbl2_hscr_n_243);
  lbl2_hscr_g18772 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_195, A2 => lbl2_hscr_n_116, A3 => lbl2_hscr_n_13, ZN => lbl2_hscr_n_242);
  lbl2_hscr_g18773 : CKND1BWP7T port map(I => lbl2_hscr_n_0, ZN => lbl2_hscr_n_237);
  lbl2_hscr_g18774 : INVD1BWP7T port map(I => lbl2_hscr_n_228, ZN => lbl2_hscr_n_227);
  lbl2_hscr_g18775 : OAI221D0BWP7T port map(A1 => lbl2_hscr_n_158, A2 => lbl2_hscr_n_64, B1 => lbl2_v_count(0), B2 => lbl2_hscr_n_99, C => lbl2_hscr_n_117, ZN => lbl2_hscr_n_225);
  lbl2_hscr_g18776 : NR2D0BWP7T port map(A1 => lbl2_hscr_n_193, A2 => lbl2_hscr_n_123, ZN => lbl2_hscr_n_224);
  lbl2_hscr_g18778 : AN2D0BWP7T port map(A1 => lbl2_hscr_n_205, A2 => lbl2_hscr_n_171, Z => lbl2_hscr_n_236);
  lbl2_hscr_g18779 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_117, B1 => lbl2_hscr_n_194, ZN => lbl2_hscr_n_235);
  lbl2_hscr_g18780 : NR2D0BWP7T port map(A1 => lbl2_hscr_n_193, A2 => lbl2_hscr_n_139, ZN => lbl2_hscr_n_234);
  lbl2_hscr_g18781 : OR2D1BWP7T port map(A1 => lbl2_hscr_n_197, A2 => lbl2_hscr_n_68, Z => lbl2_hscr_n_233);
  lbl2_hscr_g18782 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_193, A2 => lbl2_hscr_n_68, ZN => lbl2_hscr_n_232);
  lbl2_hscr_g18783 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_194, A2 => lbl2_v_count(0), ZN => lbl2_hscr_n_231);
  lbl2_hscr_g18784 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_194, A2 => lbl2_hscr_n_64, ZN => lbl2_hscr_n_230);
  lbl2_hscr_g18785 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_194, A2 => lbl2_v_count(1), ZN => lbl2_hscr_n_229);
  lbl2_hscr_g18786 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_194, A2 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_228);
  lbl2_hscr_g18787 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_196, A2 => lbl2_hscr_n_145, ZN => lbl2_hscr_n_226);
  lbl2_hscr_g18788 : OAI211D1BWP7T port map(A1 => lbl2_h_count(3), A2 => lbl2_hscr_n_45, B => lbl2_hscr_n_179, C => lbl2_hscr_n_88, ZN => lbl2_hscr_n_219);
  lbl2_hscr_g18789 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_80, A2 => lbl2_hscr_n_55, B => lbl2_hscr_n_194, ZN => lbl2_hscr_n_218);
  lbl2_hscr_g18790 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_76, A2 => lbl2_hscr_n_80, B => lbl2_hscr_n_204, ZN => lbl2_hscr_n_217);
  lbl2_hscr_g18791 : AO21D0BWP7T port map(A1 => lbl2_hscr_n_172, A2 => lbl2_hscr_n_80, B => lbl2_hscr_n_108, Z => lbl2_hscr_n_216);
  lbl2_hscr_g18792 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_133, A2 => lbl2_hscr_n_118, B => lbl2_hscr_n_202, ZN => lbl2_hscr_n_215);
  lbl2_hscr_g18793 : OR3XD1BWP7T port map(A1 => lbl2_hscr_n_104, A2 => lbl2_hscr_n_155, A3 => lbl2_hscr_n_193, Z => lbl2_hscr_n_214);
  lbl2_hscr_g18794 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_104, B1 => lbl2_hscr_n_172, B2 => lbl2_hscr_n_183, ZN => lbl2_hscr_n_213);
  lbl2_hscr_g18795 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_176, A2 => lbl2_hscr_n_162, B => lbl2_hscr_n_199, ZN => lbl2_hscr_n_212);
  lbl2_hscr_g18796 : AO21D0BWP7T port map(A1 => lbl2_hscr_n_158, A2 => lbl2_hscr_n_142, B => lbl2_hscr_n_207, Z => lbl2_hscr_n_211);
  lbl2_hscr_g18797 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_182, A2 => lbl2_hscr_n_120, A3 => lbl2_hscr_n_67, ZN => lbl2_hscr_n_223);
  lbl2_hscr_g18798 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_120, A2 => lbl2_hscr_n_98, B => lbl2_hscr_n_194, ZN => lbl2_hscr_n_222);
  lbl2_hscr_g18799 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_180, A2 => lbl2_hscr_n_132, A3 => lbl2_hscr_n_172, ZN => lbl2_hscr_n_221);
  lbl2_hscr_g18800 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_173, B1 => lbl2_hscr_n_82, B2 => lbl2_hscr_n_116, ZN => lbl2_hscr_n_220);
  lbl2_hscr_g18801 : INVD1BWP7T port map(I => lbl2_hscr_n_201, ZN => lbl2_hscr_n_202);
  lbl2_hscr_g18802 : INVD1BWP7T port map(I => lbl2_hscr_n_200, ZN => lbl2_hscr_n_199);
  lbl2_hscr_g18803 : INR2D1BWP7T port map(A1 => lbl2_hscr_n_183, B1 => lbl2_hscr_n_138, ZN => lbl2_hscr_n_210);
  lbl2_hscr_g18804 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_186, A2 => lbl2_h_count(2), ZN => lbl2_hscr_n_209);
  lbl2_hscr_g18805 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_182, A2 => FE_DBTN20_lbl2_h_count_2, ZN => lbl2_hscr_n_208);
  lbl2_hscr_g18806 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_186, A2 => FE_DBTN20_lbl2_h_count_2, ZN => lbl2_hscr_n_207);
  lbl2_hscr_g18807 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_175, A2 => lbl2_hscr_n_159, ZN => lbl2_hscr_n_206);
  lbl2_hscr_g18808 : INR2D1BWP7T port map(A1 => lbl2_hscr_n_180, B1 => lbl2_hscr_n_132, ZN => lbl2_hscr_n_205);
  lbl2_hscr_g18809 : AN2D1BWP7T port map(A1 => lbl2_hscr_n_180, A2 => lbl2_hscr_n_132, Z => lbl2_hscr_n_204);
  lbl2_hscr_g18810 : INR2XD0BWP7T port map(A1 => lbl2_hscr_n_92, B1 => lbl2_hscr_n_185, ZN => lbl2_hscr_n_203);
  lbl2_hscr_g18811 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_160, A2 => lbl2_hscr_n_172, ZN => lbl2_hscr_n_201);
  lbl2_hscr_g18812 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_183, A2 => lbl2_hscr_n_103, ZN => lbl2_hscr_n_200);
  lbl2_hscr_g18814 : INVD1BWP7T port map(I => lbl2_hscr_n_194, ZN => lbl2_hscr_n_193);
  lbl2_hscr_g18815 : AO31D1BWP7T port map(A1 => lbl2_hscr_n_145, A2 => lbl2_hscr_n_76, A3 => lbl2_hscr_n_48, B => lbl2_hscr_n_165, Z => lbl2_hscr_n_192);
  lbl2_hscr_g18816 : MOAI22D0BWP7T port map(A1 => lbl2_hscr_n_132, A2 => lbl2_hscr_n_134, B1 => lbl2_hscr_n_146, B2 => lbl2_hscr_n_160, ZN => lbl2_hscr_n_191);
  lbl2_hscr_g18817 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_161, B1 => lbl2_hscr_n_118, B2 => lbl2_hscr_n_160, ZN => lbl2_hscr_n_190);
  lbl2_hscr_g18818 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_39, A2 => lbl2_hscr_n_27, A3 => lbl2_v_count(2), B => lbl2_hscr_n_166, ZN => lbl2_hscr_n_189);
  lbl2_hscr_g18819 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_157, A2 => lbl2_hscr_n_98, B => FE_DBTN20_lbl2_h_count_2, ZN => lbl2_hscr_n_188);
  lbl2_hscr_g18820 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_99, A2 => lbl2_hscr_n_46, B => lbl2_hscr_n_181, ZN => lbl2_hscr_n_187);
  lbl2_hscr_g18821 : NR2D0BWP7T port map(A1 => lbl2_hscr_n_171, A2 => lbl2_hscr_n_64, ZN => lbl2_hscr_n_198);
  lbl2_hscr_g18822 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_135, B1 => lbl2_hscr_n_172, B2 => lbl2_hscr_n_153, ZN => lbl2_hscr_n_197);
  lbl2_hscr_g18823 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_132, A2 => lbl2_hscr_n_171, ZN => lbl2_hscr_n_196);
  lbl2_hscr_g18824 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_131, A2 => lbl2_hscr_n_171, A3 => lbl2_hscr_n_104, ZN => lbl2_hscr_n_195);
  lbl2_hscr_g18825 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_131, A2 => lbl2_hscr_n_172, ZN => lbl2_hscr_n_194);
  lbl2_hscr_g18826 : INVD0BWP7T port map(I => lbl2_hscr_n_182, ZN => lbl2_hscr_n_181);
  lbl2_hscr_g18827 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_70, A2 => lbl2_hscr_n_19, A3 => lbl2_hscr_n_9, B => lbl2_hscr_n_400, ZN => lbl2_hscr_n_179);
  lbl2_hscr_g18828 : OR2D1BWP7T port map(A1 => lbl2_hscr_n_162, A2 => lbl2_hscr_n_120, Z => lbl2_hscr_n_178);
  lbl2_hscr_g18829 : IND3D1BWP7T port map(A1 => lbl2_central_x_vec(7), B1 => lbl2_hscr_n_29, B2 => lbl2_hscr_n_136, ZN => lbl2_hscr_n_177);
  lbl2_hscr_g18830 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_154, A2 => lbl2_hscr_n_101, ZN => lbl2_hscr_n_186);
  lbl2_hscr_g18831 : OAI211D1BWP7T port map(A1 => lbl2_n_123, A2 => lbl2_hscr_n_63, B => lbl2_hscr_n_136, C => lbl2_hscr_n_32, ZN => lbl2_hscr_n_185);
  lbl2_hscr_g18832 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_157, A2 => lbl2_hscr_n_131, ZN => lbl2_hscr_n_184);
  lbl2_hscr_g18833 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_154, A2 => lbl2_hscr_n_48, ZN => lbl2_hscr_n_183);
  lbl2_hscr_g18834 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_154, A2 => lbl2_hscr_n_82, ZN => lbl2_hscr_n_182);
  lbl2_hscr_g18835 : AOI211XD0BWP7T port map(A1 => lbl2_hscr_n_105, A2 => lbl2_central_x_vec(8), B => lbl2_hscr_n_129, C => lbl2_hscr_n_31, ZN => lbl2_hscr_n_180);
  lbl2_hscr_g18836 : INVD0BWP7T port map(I => lbl2_hscr_n_175, ZN => lbl2_hscr_n_174);
  lbl2_hscr_g18837 : INVD1BWP7T port map(I => lbl2_hscr_n_172, ZN => lbl2_hscr_n_171);
  lbl2_hscr_g18838 : MAOI22D0BWP7T port map(A1 => lbl2_hscr_n_47, A2 => lbl2_hscr_n_53, B1 => lbl2_hscr_n_143, B2 => lbl2_hscr_n_64, ZN => lbl2_hscr_n_170);
  lbl2_hscr_g18839 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_117, A2 => lbl2_v_count(1), B => lbl2_hscr_n_158, ZN => lbl2_hscr_n_169);
  lbl2_hscr_g18840 : AO21D0BWP7T port map(A1 => lbl2_hscr_n_133, A2 => lbl2_hscr_n_82, B => lbl2_hscr_n_163, Z => lbl2_hscr_n_168);
  lbl2_hscr_g18841 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_138, A2 => lbl2_hscr_n_2, B => lbl2_hscr_n_164, ZN => lbl2_hscr_n_167);
  lbl2_hscr_g18842 : OAI211D1BWP7T port map(A1 => lbl2_hscr_n_39, A2 => lbl2_hscr_n_130, B => lbl2_hscr_n_113, C => lbl2_hscr_n_112, ZN => lbl2_hscr_n_166);
  lbl2_hscr_g18843 : MOAI22D0BWP7T port map(A1 => lbl2_hscr_n_115, A2 => lbl2_hscr_n_145, B1 => lbl2_hscr_n_100, B2 => lbl2_hscr_n_50, ZN => lbl2_hscr_n_165);
  lbl2_hscr_g18844 : MOAI22D0BWP7T port map(A1 => lbl2_hscr_n_139, A2 => lbl2_hscr_n_2, B1 => lbl2_hscr_n_120, B2 => lbl2_hscr_n_13, ZN => lbl2_hscr_n_176);
  lbl2_hscr_g18845 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_131, A2 => lbl2_hscr_n_139, A3 => lbl2_v_count(0), ZN => lbl2_hscr_n_175);
  lbl2_hscr_g18846 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_133, A2 => lbl2_hscr_n_132, A3 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_173);
  lbl2_hscr_g18847 : MOAI22D1BWP7T port map(A1 => lbl2_hscr_n_109, A2 => lbl2_central_x_vec(6), B1 => lbl2_hscr_n_109, B2 => lbl2_central_x_vec(6), ZN => lbl2_hscr_n_172);
  lbl2_hscr_g18848 : INVD1BWP7T port map(I => lbl2_hscr_n_158, ZN => lbl2_hscr_n_157);
  lbl2_hscr_g18849 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_137, A2 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_164);
  lbl2_hscr_g18850 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_141, A2 => lbl2_v_count(1), ZN => lbl2_hscr_n_163);
  lbl2_hscr_g18851 : AN2D0BWP7T port map(A1 => lbl2_hscr_n_137, A2 => lbl2_v_count(0), Z => lbl2_hscr_n_162);
  lbl2_hscr_g18852 : NR2D0BWP7T port map(A1 => lbl2_hscr_n_101, A2 => lbl2_hscr_n_145, ZN => lbl2_hscr_n_156);
  lbl2_hscr_g18853 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_145, A2 => lbl2_hscr_n_82, ZN => lbl2_hscr_n_161);
  lbl2_hscr_g18854 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_132, A2 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_160);
  lbl2_hscr_g18855 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_145, A2 => lbl2_hscr_n_82, ZN => lbl2_hscr_n_159);
  lbl2_hscr_g18856 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_140, A2 => lbl2_v_count(0), ZN => lbl2_hscr_n_158);
  lbl2_hscr_g18857 : INVD0BWP7T port map(I => lbl2_hscr_n_154, ZN => lbl2_hscr_n_153);
  lbl2_hscr_g18859 : AOI33D1BWP7T port map(A1 => lbl2_hscr_n_72, A2 => lbl2_hscr_n_23, A3 => lbl2_hscr_n_1, B1 => lbl2_hscr_n_89, B2 => lbl2_h_count(1), B3 => lbl2_h_count(3), ZN => lbl2_hscr_n_151);
  lbl2_hscr_g18860 : AOI221D0BWP7T port map(A1 => lbl2_hscr_n_60, A2 => lbl2_hscr_n_70, B1 => lbl2_hscr_n_95, B2 => lbl2_v_count(1), C => lbl2_hscr_n_128, ZN => lbl2_hscr_n_150);
  lbl2_hscr_g18861 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_123, A2 => lbl2_v_count(0), B => lbl2_hscr_n_53, ZN => lbl2_hscr_n_149);
  lbl2_hscr_g18862 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_107, A2 => lbl2_hscr_n_13, B => lbl2_hscr_n_144, ZN => lbl2_hscr_n_148);
  lbl2_hscr_g18863 : OA21D0BWP7T port map(A1 => lbl2_hscr_n_125, A2 => lbl2_hscr_n_2, B => lbl2_hscr_n_134, Z => lbl2_hscr_n_147);
  lbl2_hscr_g18864 : OAI211D1BWP7T port map(A1 => lbl2_v_count(1), A2 => lbl2_hscr_n_99, B => lbl2_hscr_n_121, C => lbl2_hscr_n_96, ZN => lbl2_hscr_n_146);
  lbl2_hscr_g18865 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_90, B1 => lbl2_hscr_n_145, ZN => lbl2_hscr_n_155);
  lbl2_hscr_g18866 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_132, A2 => lbl2_hscr_n_116, ZN => lbl2_hscr_n_154);
  lbl2_hscr_g18867 : INVD1BWP7T port map(I => lbl2_hscr_n_116, ZN => lbl2_hscr_n_145);
  lbl2_hscr_g18868 : INR2D1BWP7T port map(A1 => lbl2_hscr_n_118, B1 => lbl2_hscr_n_13, ZN => lbl2_hscr_n_144);
  lbl2_hscr_g18869 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_120, A2 => lbl2_hscr_n_1, ZN => lbl2_hscr_n_143);
  lbl2_hscr_g18870 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_122, A2 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_142);
  lbl2_hscr_g18871 : OR2D1BWP7T port map(A1 => lbl2_hscr_n_117, A2 => lbl2_hscr_n_2, Z => lbl2_hscr_n_141);
  lbl2_hscr_g18872 : AN2D1BWP7T port map(A1 => lbl2_hscr_n_118, A2 => lbl2_hscr_n_1, Z => lbl2_hscr_n_140);
  lbl2_hscr_g18873 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_118, A2 => lbl2_v_count(1), ZN => lbl2_hscr_n_139);
  lbl2_hscr_g18874 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_122, A2 => lbl2_v_count(1), ZN => lbl2_hscr_n_138);
  lbl2_hscr_g18875 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_121, A2 => lbl2_v_count(1), ZN => lbl2_hscr_n_137);
  lbl2_hscr_g18876 : INVD1BWP7T port map(I => lbl2_hscr_n_134, ZN => lbl2_hscr_n_133);
  lbl2_hscr_g18877 : INVD1BWP7T port map(I => lbl2_hscr_n_132, ZN => lbl2_hscr_n_131);
  lbl2_hscr_g18878 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_86, A2 => lbl2_h_count(3), B1 => lbl2_hscr_n_27, B2 => FE_DBTN18_lbl2_v_count_2, ZN => lbl2_hscr_n_130);
  lbl2_hscr_g18879 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_105, A2 => lbl2_central_x_vec(8), A3 => lbl2_central_x_vec(7), ZN => lbl2_hscr_n_129);
  lbl2_hscr_g18880 : OAI33D1BWP7T port map(A1 => lbl2_v_count(0), A2 => lbl2_hscr_n_33, A3 => lbl2_hscr_n_81, B1 => lbl2_v_count(2), B2 => lbl2_hscr_n_36, B3 => lbl2_hscr_n_74, ZN => lbl2_hscr_n_128);
  lbl2_hscr_g18881 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_97, A2 => lbl2_v_count(1), B => lbl2_hscr_n_120, ZN => lbl2_hscr_n_127);
  lbl2_hscr_g18882 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_77, A2 => lbl2_hscr_n_17, A3 => lbl2_h_count(1), B1 => lbl2_hscr_n_85, B2 => lbl2_hscr_n_29, ZN => lbl2_hscr_n_126);
  lbl2_hscr_g18883 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_87, A2 => lbl2_hscr_n_78, A3 => lbl2_hscr_n_35, ZN => lbl2_hscr_n_136);
  lbl2_hscr_g18884 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_104, B1 => lbl2_hscr_n_1, B2 => lbl2_hscr_n_65, ZN => lbl2_hscr_n_135);
  lbl2_hscr_g18885 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_107, A2 => lbl2_hscr_n_83, A3 => lbl2_v_count(1), ZN => lbl2_hscr_n_134);
  lbl2_hscr_g18886 : MOAI22D0BWP7T port map(A1 => lbl2_hscr_n_105, A2 => lbl2_central_x_vec(7), B1 => lbl2_hscr_n_105, B2 => lbl2_central_x_vec(7), ZN => lbl2_hscr_n_132);
  lbl2_hscr_g18887 : INVD1BWP7T port map(I => lbl2_hscr_n_122, ZN => lbl2_hscr_n_121);
  lbl2_hscr_g18888 : INVD1BWP7T port map(I => lbl2_hscr_n_119, ZN => lbl2_hscr_n_120);
  lbl2_hscr_g18889 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_98, A2 => lbl2_hscr_n_97, ZN => lbl2_hscr_n_125);
  lbl2_hscr_g18890 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_97, A2 => lbl2_hscr_n_48, ZN => lbl2_hscr_n_124);
  lbl2_hscr_g18891 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_98, A2 => lbl2_v_count(1), ZN => lbl2_hscr_n_123);
  lbl2_hscr_g18892 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_99, A2 => lbl2_hscr_n_41, ZN => lbl2_hscr_n_122);
  lbl2_hscr_g18893 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_97, A2 => lbl2_hscr_n_41, ZN => lbl2_hscr_n_119);
  lbl2_hscr_g18894 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_96, A2 => lbl2_hscr_n_41, ZN => lbl2_hscr_n_118);
  lbl2_hscr_g18895 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_98, A2 => lbl2_hscr_n_41, ZN => lbl2_hscr_n_117);
  lbl2_hscr_g18896 : AOI31D0BWP7T port map(A1 => lbl2_hscr_n_50, A2 => lbl2_hscr_n_47, A3 => lbl2_v_count(3), B => lbl2_hscr_n_25, ZN => lbl2_hscr_n_115);
  lbl2_hscr_g18897 : AO21D0BWP7T port map(A1 => lbl2_hscr_n_82, A2 => lbl2_hscr_n_50, B => lbl2_hscr_n_54, Z => lbl2_hscr_n_114);
  lbl2_hscr_g18898 : OAI211D1BWP7T port map(A1 => FE_DBTN18_lbl2_v_count_2, A2 => lbl2_hscr_n_15, B => lbl2_hscr_n_77, C => lbl2_h_count(1), ZN => lbl2_hscr_n_113);
  lbl2_hscr_g18899 : IND4D0BWP7T port map(A1 => lbl2_hscr_n_62, B1 => lbl2_v_count(1), B2 => lbl2_hscr_n_14, B3 => lbl2_hscr_n_40, ZN => lbl2_hscr_n_112);
  lbl2_hscr_g18900 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_34, A2 => lbl2_hscr_n_13, A3 => lbl2_hscr_n_15, B1 => lbl2_hscr_n_401, B2 => lbl2_hscr_n_18, ZN => lbl2_hscr_n_111);
  lbl2_hscr_g18901 : OAI31D0BWP7T port map(A1 => lbl2_v_count(6), A2 => lbl2_v_count(2), A3 => lbl2_hscr_n_12, B => lbl2_hscr_n_93, ZN => lbl2_hscr_n_110);
  lbl2_hscr_g18902 : MAOI22D1BWP7T port map(A1 => lbl2_hscr_n_49, A2 => lbl2_central_x_vec(5), B1 => lbl2_hscr_n_49, B2 => lbl2_central_x_vec(5), ZN => lbl2_hscr_n_116);
  lbl2_hscr_g18903 : INVD0BWP7T port map(I => lbl2_hscr_n_107, ZN => lbl2_hscr_n_106);
  lbl2_hscr_g18904 : INVD0BWP7T port map(I => lbl2_hscr_n_103, ZN => lbl2_hscr_n_102);
  lbl2_hscr_g18905 : INVD0BWP7T port map(I => lbl2_hscr_n_101, ZN => lbl2_hscr_n_100);
  lbl2_hscr_g18906 : INVD1BWP7T port map(I => lbl2_hscr_n_99, ZN => lbl2_hscr_n_98);
  lbl2_hscr_g18907 : INVD1BWP7T port map(I => lbl2_hscr_n_97, ZN => lbl2_hscr_n_96);
  lbl2_hscr_g18908 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_49, B1 => lbl2_central_x_vec(5), ZN => lbl2_hscr_n_109);
  lbl2_hscr_g18909 : AN2D1BWP7T port map(A1 => lbl2_hscr_n_76, A2 => lbl2_v_count(3), Z => lbl2_hscr_n_108);
  lbl2_hscr_g18910 : INR2D1BWP7T port map(A1 => lbl2_hscr_n_41, B1 => lbl2_hscr_n_79, ZN => lbl2_hscr_n_107);
  lbl2_hscr_g18911 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_22, A2 => lbl2_hscr_n_49, ZN => lbl2_hscr_n_105);
  lbl2_hscr_g18912 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_41, B1 => lbl2_hscr_n_79, ZN => lbl2_hscr_n_104);
  lbl2_hscr_g18913 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_64, A2 => lbl2_h_count(2), ZN => lbl2_hscr_n_103);
  lbl2_hscr_g18914 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_64, A2 => lbl2_hscr_n_48, ZN => lbl2_hscr_n_101);
  lbl2_hscr_g18915 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_79, A2 => lbl2_hscr_n_83, ZN => lbl2_hscr_n_99);
  lbl2_hscr_g18916 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_79, A2 => lbl2_hscr_n_83, ZN => lbl2_hscr_n_97);
  lbl2_hscr_g18917 : INVD0BWP7T port map(I => lbl2_hscr_n_94, ZN => lbl2_hscr_n_95);
  lbl2_hscr_g18918 : CKND1BWP7T port map(I => lbl2_hscr_n_92, ZN => lbl2_hscr_n_93);
  lbl2_hscr_g18919 : MOAI22D0BWP7T port map(A1 => lbl2_hscr_n_14, A2 => lbl2_hscr_n_1, B1 => lbl2_hscr_n_39, B2 => lbl2_hscr_n_18, ZN => lbl2_hscr_n_89);
  lbl2_hscr_g18920 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_70, A2 => lbl2_hscr_n_42, B1 => lbl2_hscr_n_61, B2 => lbl2_hscr_n_29, ZN => lbl2_hscr_n_88);
  lbl2_hscr_g18921 : AOI211XD0BWP7T port map(A1 => lbl2_hscr_n_44, A2 => lbl2_h_count(3), B => lbl2_central_x_vec(8), C => lbl2_central_x_vec(7), ZN => lbl2_hscr_n_87);
  lbl2_hscr_g18922 : OAI31D0BWP7T port map(A1 => FE_DBTN19_lbl2_h_count_1, A2 => FE_DBTN18_lbl2_v_count_2, A3 => lbl2_hscr_n_43, B => lbl2_hscr_n_14, ZN => lbl2_hscr_n_86);
  lbl2_hscr_g18923 : IOA21D0BWP7T port map(A1 => lbl2_hscr_n_18, A2 => lbl2_v_count(0), B => lbl2_hscr_n_45, ZN => lbl2_hscr_n_85);
  lbl2_hscr_g18924 : AOI32D1BWP7T port map(A1 => lbl2_hscr_n_11, A2 => lbl2_hscr_n_37, A3 => lbl2_h_count(1), B1 => lbl2_hscr_n_70, B2 => lbl2_hscr_n_13, ZN => lbl2_hscr_n_84);
  lbl2_hscr_g18925 : IND3D1BWP7T port map(A1 => lbl2_hscr_n_21, B1 => lbl2_v_count(0), B2 => lbl2_hscr_n_72, ZN => lbl2_hscr_n_94);
  lbl2_hscr_g18926 : ND3D0BWP7T port map(A1 => lbl2_hscr_n_73, A2 => lbl2_v_count(7), A3 => lbl2_v_count(8), ZN => lbl2_hscr_n_92);
  lbl2_hscr_g18927 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_64, A2 => lbl2_hscr_n_47, ZN => lbl2_hscr_n_91);
  lbl2_hscr_g18928 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_82, A2 => lbl2_hscr_n_48, ZN => lbl2_hscr_n_90);
  lbl2_hscr_g18929 : INVD1BWP7T port map(I => lbl2_hscr_n_65, ZN => lbl2_hscr_n_83);
  lbl2_hscr_g18930 : INVD1BWP7T port map(I => lbl2_hscr_n_64, ZN => lbl2_hscr_n_82);
  lbl2_hscr_g18931 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_54, A2 => lbl2_hscr_n_10, B => lbl2_v_count(8), ZN => lbl2_hscr_n_78);
  lbl2_hscr_g18932 : IND2D1BWP7T port map(A1 => lbl2_hscr_n_42, B1 => lbl2_hscr_n_72, ZN => lbl2_hscr_n_81);
  lbl2_hscr_g18933 : INR2D1BWP7T port map(A1 => lbl2_hscr_n_50, B1 => lbl2_v_count(3), ZN => lbl2_hscr_n_80);
  lbl2_hscr_g18934 : OA211D0BWP7T port map(A1 => lbl2_v_count(4), A2 => lbl2_hscr_n_17, B => lbl2_hscr_n_46, C => lbl2_hscr_n_30, Z => lbl2_hscr_n_79);
  lbl2_hscr_g18936 : OA21D0BWP7T port map(A1 => lbl2_hscr_n_43, A2 => FE_DBTN19_lbl2_h_count_1, B => lbl2_hscr_n_40, Z => lbl2_hscr_n_74);
  lbl2_hscr_g18937 : NR3D0BWP7T port map(A1 => lbl2_hscr_n_40, A2 => lbl2_hscr_n_21, A3 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_77);
  lbl2_hscr_g18938 : AN3D1BWP7T port map(A1 => lbl2_hscr_n_50, A2 => lbl2_hscr_n_30, A3 => lbl2_hscr_n_26, Z => lbl2_hscr_n_76);
  lbl2_hscr_g18939 : INVD0BWP7T port map(I => lbl2_hscr_n_68, ZN => lbl2_hscr_n_67);
  lbl2_hscr_g18940 : AOI211D1BWP7T port map(A1 => lbl2_central_x_vec(5), A2 => lbl2_h_count(4), B => lbl2_hscr_n_20, C => lbl2_hscr_n_24, ZN => lbl2_hscr_n_66);
  lbl2_hscr_g18941 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_52, A2 => lbl2_hscr_n_10, ZN => lbl2_hscr_n_73);
  lbl2_hscr_g18942 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_56, A2 => lbl2_hscr_n_40, ZN => lbl2_hscr_n_72);
  lbl2_hscr_g18943 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_48, A2 => lbl2_h_count(2), ZN => lbl2_hscr_n_71);
  lbl2_hscr_g18944 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_57, A2 => lbl2_hscr_n_39, ZN => lbl2_hscr_n_70);
  lbl2_hscr_g18946 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_47, A2 => lbl2_h_count(2), ZN => lbl2_hscr_n_68);
  lbl2_hscr_g18947 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_22, A2 => FE_DBTN21_lbl2_h_count_3, B => lbl2_hscr_n_44, ZN => lbl2_hscr_n_63);
  lbl2_hscr_g18948 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_34, A2 => lbl2_v_count(0), B => lbl2_hscr_n_23, ZN => lbl2_hscr_n_62);
  lbl2_hscr_g18949 : MOAI22D0BWP7T port map(A1 => lbl2_hscr_n_12, A2 => lbl2_h_count(3), B1 => lbl2_hscr_n_19, B2 => lbl2_v_count(1), ZN => lbl2_hscr_n_61);
  lbl2_hscr_g18950 : MOAI22D0BWP7T port map(A1 => lbl2_hscr_n_12, A2 => lbl2_hscr_n_21, B1 => lbl2_hscr_n_29, B2 => lbl2_hscr_n_19, ZN => lbl2_hscr_n_60);
  lbl2_hscr_g18951 : IAO21D0BWP7T port map(A1 => lbl2_hscr_n_35, A2 => lbl2_v_count(5), B => lbl2_v_count(4), ZN => lbl2_hscr_n_59);
  lbl2_hscr_g18952 : MOAI22D0BWP7T port map(A1 => lbl2_central_x_vec(7), A2 => lbl2_hscr_n_20, B1 => lbl2_central_x_vec(6), B2 => lbl2_hscr_n_20, ZN => lbl2_hscr_n_58);
  lbl2_hscr_g18953 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_16, A2 => lbl2_v_count(3), B => lbl2_hscr_n_53, ZN => lbl2_hscr_n_65);
  lbl2_hscr_g18954 : AOI21D1BWP7T port map(A1 => lbl2_hscr_n_28, A2 => lbl2_h_count(4), B => lbl2_hscr_n_49, ZN => lbl2_hscr_n_64);
  lbl2_hscr_g18955 : INVD0BWP7T port map(I => lbl2_hscr_n_56, ZN => lbl2_hscr_n_57);
  lbl2_hscr_g18956 : INVD1BWP7T port map(I => lbl2_hscr_n_52, ZN => lbl2_hscr_n_51);
  lbl2_hscr_g18957 : INVD1BWP7T port map(I => lbl2_hscr_n_48, ZN => lbl2_hscr_n_47);
  lbl2_hscr_g18958 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_37, A2 => lbl2_hscr_n_15, ZN => lbl2_hscr_n_56);
  lbl2_hscr_g18959 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_26, A2 => lbl2_v_count(5), ZN => lbl2_hscr_n_55);
  lbl2_hscr_g18960 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_30, A2 => lbl2_v_count(5), ZN => lbl2_hscr_n_54);
  lbl2_hscr_g18961 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_16, A2 => lbl2_v_count(3), ZN => lbl2_hscr_n_53);
  lbl2_hscr_g18962 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_25, A2 => lbl2_v_count(5), ZN => lbl2_hscr_n_52);
  lbl2_hscr_g18963 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_26, A2 => lbl2_v_count(5), ZN => lbl2_hscr_n_50);
  lbl2_hscr_g18964 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_28, A2 => lbl2_h_count(4), ZN => lbl2_hscr_n_49);
  lbl2_hscr_g18965 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_28, A2 => lbl2_hscr_n_36, ZN => lbl2_hscr_n_48);
  lbl2_hscr_g18966 : INVD1BWP7T port map(I => lbl2_hscr_n_40, ZN => lbl2_hscr_n_39);
  lbl2_hscr_g18968 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_17, A2 => lbl2_hscr_n_25, ZN => lbl2_hscr_n_46);
  lbl2_hscr_g18969 : CKND2D0BWP7T port map(A1 => lbl2_hscr_n_11, A2 => lbl2_v_count(2), ZN => lbl2_hscr_n_45);
  lbl2_hscr_g18970 : INR2D1BWP7T port map(A1 => lbl2_h_count(4), B1 => lbl2_hscr_n_22, ZN => lbl2_hscr_n_44);
  lbl2_hscr_g18971 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_2, A2 => lbl2_h_count(0), B => lbl2_hscr_n_1, ZN => lbl2_hscr_n_43);
  lbl2_hscr_g18972 : AOI22D0BWP7T port map(A1 => lbl2_hscr_n_1, A2 => lbl2_h_count(1), B1 => lbl2_v_count(1), B2 => FE_DBTN19_lbl2_h_count_1, ZN => lbl2_hscr_n_42);
  lbl2_hscr_g18973 : AOI21D0BWP7T port map(A1 => lbl2_hscr_n_1, A2 => lbl2_v_count(2), B => lbl2_hscr_n_18, ZN => lbl2_hscr_n_41);
  lbl2_hscr_g18974 : MAOI22D0BWP7T port map(A1 => lbl2_v_count(2), A2 => lbl2_v_count(3), B1 => lbl2_v_count(2), B2 => lbl2_v_count(3), ZN => lbl2_hscr_n_40);
  lbl2_hscr_g18975 : INVD0BWP7T port map(I => lbl2_hscr_n_34, ZN => lbl2_hscr_n_33);
  lbl2_hscr_g18976 : INVD0BWP7T port map(I => lbl2_hscr_n_32, ZN => lbl2_hscr_n_31);
  lbl2_hscr_g18977 : INVD0BWP7T port map(I => lbl2_hscr_n_28, ZN => lbl2_hscr_n_27);
  lbl2_hscr_g18978 : INVD1BWP7T port map(I => lbl2_hscr_n_26, ZN => lbl2_hscr_n_25);
  lbl2_hscr_g18979 : NR2XD0BWP7T port map(A1 => lbl2_h_count(4), A2 => direction_between(2), ZN => lbl2_hscr_n_24);
  lbl2_hscr_g18980 : NR2D0BWP7T port map(A1 => lbl2_h_count(2), A2 => lbl2_v_count(2), ZN => lbl2_hscr_n_37);
  lbl2_hscr_g18981 : ND2D1BWP7T port map(A1 => lbl2_h_count(2), A2 => lbl2_h_count(3), ZN => lbl2_hscr_n_36);
  lbl2_hscr_g18982 : NR2XD0BWP7T port map(A1 => lbl2_v_count(7), A2 => lbl2_v_count(8), ZN => lbl2_hscr_n_35);
  lbl2_hscr_g18983 : NR2D0BWP7T port map(A1 => lbl2_h_count(3), A2 => lbl2_h_count(0), ZN => lbl2_hscr_n_34);
  lbl2_hscr_g18984 : ND2D1BWP7T port map(A1 => lbl2_central_x_vec(8), A2 => lbl2_central_x_vec(7), ZN => lbl2_hscr_n_32);
  lbl2_hscr_g18985 : OR2D1BWP7T port map(A1 => lbl2_v_count(3), A2 => lbl2_v_count(4), Z => lbl2_hscr_n_30);
  lbl2_hscr_g18986 : NR2D1BWP7T port map(A1 => lbl2_h_count(1), A2 => lbl2_h_count(0), ZN => lbl2_hscr_n_29);
  lbl2_hscr_g18987 : CKND2D1BWP7T port map(A1 => FE_DBTN21_lbl2_h_count_3, A2 => FE_DBTN20_lbl2_h_count_2, ZN => lbl2_hscr_n_28);
  lbl2_hscr_g18988 : CKND2D1BWP7T port map(A1 => lbl2_v_count(4), A2 => lbl2_v_count(3), ZN => lbl2_hscr_n_26);
  lbl2_hscr_g18989 : INVD0BWP7T port map(I => lbl2_hscr_n_17, ZN => lbl2_hscr_n_16);
  lbl2_hscr_g18990 : INVD0BWP7T port map(I => lbl2_hscr_n_15, ZN => lbl2_hscr_n_14);
  lbl2_hscr_g18991 : INVD0BWP7T port map(I => lbl2_hscr_n_12, ZN => lbl2_hscr_n_11);
  lbl2_hscr_g18992 : NR2D0BWP7T port map(A1 => lbl2_h_count(3), A2 => lbl2_h_count(1), ZN => lbl2_hscr_n_23);
  lbl2_hscr_g18993 : ND2D1BWP7T port map(A1 => lbl2_central_x_vec(6), A2 => lbl2_central_x_vec(5), ZN => lbl2_hscr_n_22);
  lbl2_hscr_g18994 : ND2D1BWP7T port map(A1 => lbl2_h_count(3), A2 => lbl2_h_count(0), ZN => lbl2_hscr_n_21);
  lbl2_hscr_g18995 : NR2XD0BWP7T port map(A1 => lbl2_central_x_vec(5), A2 => lbl2_h_count(4), ZN => lbl2_hscr_n_20);
  lbl2_hscr_g18996 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_2, A2 => lbl2_h_count(3), ZN => lbl2_hscr_n_19);
  lbl2_hscr_g18997 : NR2D1BWP7T port map(A1 => lbl2_hscr_n_1, A2 => lbl2_v_count(2), ZN => lbl2_hscr_n_18);
  lbl2_hscr_g18998 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_1, A2 => FE_DBTN18_lbl2_v_count_2, ZN => lbl2_hscr_n_17);
  lbl2_hscr_g18999 : NR2D1BWP7T port map(A1 => FE_DBTN20_lbl2_h_count_2, A2 => FE_DBTN18_lbl2_v_count_2, ZN => lbl2_hscr_n_15);
  lbl2_hscr_g19000 : NR2XD0BWP7T port map(A1 => lbl2_hscr_n_1, A2 => lbl2_v_count(0), ZN => lbl2_hscr_n_13);
  lbl2_hscr_g19001 : ND2D1BWP7T port map(A1 => lbl2_hscr_n_1, A2 => lbl2_hscr_n_2, ZN => lbl2_hscr_n_12);
  lbl2_hscr_g19002 : INVD1BWP7T port map(I => lbl2_v_count(6), ZN => lbl2_hscr_n_10);
  lbl2_hscr_g19003 : INVD1BWP7T port map(I => lbl2_h_count(0), ZN => lbl2_hscr_n_9);
  lbl2_hscr_g19006 : INVD0BWP7T port map(I => lbl2_central_x_vec(6), ZN => lbl2_hscr_n_6);
  lbl2_hscr_g19010 : INVD1BWP7T port map(I => lbl2_v_count(0), ZN => lbl2_hscr_n_2);
  lbl2_hscr_g19011 : INVD1BWP7T port map(I => lbl2_v_count(1), ZN => lbl2_hscr_n_1);
  lbl2_hscr_g2 : INR2D1BWP7T port map(A1 => lbl2_hscr_n_196, B1 => lbl2_hscr_n_139, ZN => lbl2_hscr_n_0);
  lbl2_hscr_g19012 : INVD0BWP7T port map(I => lbl2_v_count(8), ZN => lbl2_hscr_n_38);
  lbl2_hscr_g19014 : OAI21D0BWP7T port map(A1 => lbl2_hscr_n_111, A2 => lbl2_hscr_n_40, B => lbl2_hscr_n_94, ZN => lbl2_hscr_n_400);
  lbl2_hscr_g19015 : AO21D0BWP7T port map(A1 => lbl2_hscr_n_27, A2 => lbl2_hscr_n_9, B => lbl2_hscr_n_19, Z => lbl2_hscr_n_401);
  lbl5_en0_inc_add_127_23_g182 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_32, A2 => lbl5_en0_count(18), B1 => lbl5_en0_inc_add_127_23_n_32, B2 => lbl5_en0_count(18), ZN => lbl5_en0_n_298);
  lbl5_en0_inc_add_127_23_g183 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_30, A2 => lbl5_en0_count(17), B1 => lbl5_en0_inc_add_127_23_n_30, B2 => lbl5_en0_count(17), ZN => lbl5_en0_n_297);
  lbl5_en0_inc_add_127_23_g184 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_30, B1 => lbl5_en0_count(17), ZN => lbl5_en0_inc_add_127_23_n_32);
  lbl5_en0_inc_add_127_23_g185 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_28, A2 => lbl5_en0_count(16), B1 => lbl5_en0_inc_add_127_23_n_28, B2 => lbl5_en0_count(16), ZN => FE_PHN286_lbl5_en0_n_296);
  lbl5_en0_inc_add_127_23_g186 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_28, B1 => lbl5_en0_count(16), ZN => lbl5_en0_inc_add_127_23_n_30);
  lbl5_en0_inc_add_127_23_g187 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_26, A2 => lbl5_en0_count(15), B1 => lbl5_en0_inc_add_127_23_n_26, B2 => lbl5_en0_count(15), ZN => lbl5_en0_n_295);
  lbl5_en0_inc_add_127_23_g188 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_26, B1 => lbl5_en0_count(15), ZN => lbl5_en0_inc_add_127_23_n_28);
  lbl5_en0_inc_add_127_23_g189 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_24, A2 => lbl5_en0_count(14), B1 => lbl5_en0_inc_add_127_23_n_24, B2 => lbl5_en0_count(14), ZN => lbl5_en0_n_294);
  lbl5_en0_inc_add_127_23_g190 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_24, B1 => lbl5_en0_count(14), ZN => lbl5_en0_inc_add_127_23_n_26);
  lbl5_en0_inc_add_127_23_g191 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_22, A2 => lbl5_en0_count(13), B1 => lbl5_en0_inc_add_127_23_n_22, B2 => lbl5_en0_count(13), ZN => FE_PHN172_lbl5_en0_n_293);
  lbl5_en0_inc_add_127_23_g192 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_22, B1 => lbl5_en0_count(13), ZN => lbl5_en0_inc_add_127_23_n_24);
  lbl5_en0_inc_add_127_23_g193 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_20, A2 => lbl5_en0_count(12), B1 => lbl5_en0_inc_add_127_23_n_20, B2 => lbl5_en0_count(12), ZN => FE_PHN160_lbl5_en0_n_292);
  lbl5_en0_inc_add_127_23_g194 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_20, B1 => lbl5_en0_count(12), ZN => lbl5_en0_inc_add_127_23_n_22);
  lbl5_en0_inc_add_127_23_g195 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_18, A2 => lbl5_en0_count(11), B1 => lbl5_en0_inc_add_127_23_n_18, B2 => lbl5_en0_count(11), ZN => lbl5_en0_n_291);
  lbl5_en0_inc_add_127_23_g196 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_18, B1 => lbl5_en0_count(11), ZN => lbl5_en0_inc_add_127_23_n_20);
  lbl5_en0_inc_add_127_23_g197 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_16, A2 => lbl5_en0_count(10), B1 => lbl5_en0_inc_add_127_23_n_16, B2 => lbl5_en0_count(10), ZN => lbl5_en0_n_290);
  lbl5_en0_inc_add_127_23_g198 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_16, B1 => lbl5_en0_count(10), ZN => lbl5_en0_inc_add_127_23_n_18);
  lbl5_en0_inc_add_127_23_g199 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_14, A2 => lbl5_en0_count(9), B1 => lbl5_en0_inc_add_127_23_n_14, B2 => lbl5_en0_count(9), ZN => lbl5_en0_n_289);
  lbl5_en0_inc_add_127_23_g200 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_14, B1 => lbl5_en0_count(9), ZN => lbl5_en0_inc_add_127_23_n_16);
  lbl5_en0_inc_add_127_23_g201 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_12, A2 => lbl5_en0_count(8), B1 => lbl5_en0_inc_add_127_23_n_12, B2 => lbl5_en0_count(8), ZN => lbl5_en0_n_288);
  lbl5_en0_inc_add_127_23_g202 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_12, B1 => lbl5_en0_count(8), ZN => lbl5_en0_inc_add_127_23_n_14);
  lbl5_en0_inc_add_127_23_g203 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_10, A2 => lbl5_en0_count(7), B1 => lbl5_en0_inc_add_127_23_n_10, B2 => lbl5_en0_count(7), ZN => FE_PHN168_lbl5_en0_n_287);
  lbl5_en0_inc_add_127_23_g204 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_10, B1 => lbl5_en0_count(7), ZN => lbl5_en0_inc_add_127_23_n_12);
  lbl5_en0_inc_add_127_23_g205 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_8, A2 => lbl5_en0_count(6), B1 => lbl5_en0_inc_add_127_23_n_8, B2 => lbl5_en0_count(6), ZN => lbl5_en0_n_286);
  lbl5_en0_inc_add_127_23_g206 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_8, B1 => lbl5_en0_count(6), ZN => lbl5_en0_inc_add_127_23_n_10);
  lbl5_en0_inc_add_127_23_g207 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_6, A2 => lbl5_en0_count(5), B1 => lbl5_en0_inc_add_127_23_n_6, B2 => lbl5_en0_count(5), ZN => lbl5_en0_n_285);
  lbl5_en0_inc_add_127_23_g208 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_6, B1 => lbl5_en0_count(5), ZN => lbl5_en0_inc_add_127_23_n_8);
  lbl5_en0_inc_add_127_23_g209 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_4, A2 => lbl5_en0_count(4), B1 => lbl5_en0_inc_add_127_23_n_4, B2 => lbl5_en0_count(4), ZN => lbl5_en0_n_284);
  lbl5_en0_inc_add_127_23_g210 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_4, B1 => lbl5_en0_count(4), ZN => lbl5_en0_inc_add_127_23_n_6);
  lbl5_en0_inc_add_127_23_g211 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_2, A2 => lbl5_en0_count(3), B1 => lbl5_en0_inc_add_127_23_n_2, B2 => lbl5_en0_count(3), ZN => FE_PHN181_lbl5_en0_n_283);
  lbl5_en0_inc_add_127_23_g212 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_2, B1 => lbl5_en0_count(3), ZN => lbl5_en0_inc_add_127_23_n_4);
  lbl5_en0_inc_add_127_23_g213 : MOAI22D0BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_0, A2 => lbl5_en0_count(2), B1 => lbl5_en0_inc_add_127_23_n_0, B2 => lbl5_en0_count(2), ZN => lbl5_en0_n_282);
  lbl5_en0_inc_add_127_23_g214 : IND2D1BWP7T port map(A1 => lbl5_en0_inc_add_127_23_n_0, B1 => lbl5_en0_count(2), ZN => lbl5_en0_inc_add_127_23_n_2);
  lbl5_en0_inc_add_127_23_g215 : CKXOR2D0BWP7T port map(A1 => lbl5_en0_count(0), A2 => lbl5_en0_count(1), Z => lbl5_en0_n_281);
  lbl5_en0_inc_add_127_23_g216 : ND2D1BWP7T port map(A1 => lbl5_en0_count(0), A2 => lbl5_en0_count(1), ZN => lbl5_en0_inc_add_127_23_n_0);
  lbl5_en1_inc_add_127_23_g182 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_32, A2 => lbl5_en1_count(18), B1 => lbl5_en1_inc_add_127_23_n_32, B2 => lbl5_en1_count(18), ZN => FE_PHN280_lbl5_en1_n_302);
  lbl5_en1_inc_add_127_23_g183 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_30, A2 => FE_PHN185_lbl5_en1_count_17, B1 => lbl5_en1_inc_add_127_23_n_30, B2 => FE_PHN185_lbl5_en1_count_17, ZN => lbl5_en1_n_301);
  lbl5_en1_inc_add_127_23_g184 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_30, B1 => FE_PHN185_lbl5_en1_count_17, ZN => lbl5_en1_inc_add_127_23_n_32);
  lbl5_en1_inc_add_127_23_g185 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_28, A2 => FE_PHN137_lbl5_en1_count_16, B1 => lbl5_en1_inc_add_127_23_n_28, B2 => FE_PHN137_lbl5_en1_count_16, ZN => lbl5_en1_n_300);
  lbl5_en1_inc_add_127_23_g186 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_28, B1 => FE_PHN137_lbl5_en1_count_16, ZN => lbl5_en1_inc_add_127_23_n_30);
  lbl5_en1_inc_add_127_23_g187 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_26, A2 => lbl5_en1_count(15), B1 => lbl5_en1_inc_add_127_23_n_26, B2 => lbl5_en1_count(15), ZN => FE_PHN139_lbl5_en1_n_299);
  lbl5_en1_inc_add_127_23_g188 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_26, B1 => lbl5_en1_count(15), ZN => lbl5_en1_inc_add_127_23_n_28);
  lbl5_en1_inc_add_127_23_g189 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_24, A2 => lbl5_en1_count(14), B1 => lbl5_en1_inc_add_127_23_n_24, B2 => lbl5_en1_count(14), ZN => lbl5_en1_n_298);
  lbl5_en1_inc_add_127_23_g190 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_24, B1 => lbl5_en1_count(14), ZN => lbl5_en1_inc_add_127_23_n_26);
  lbl5_en1_inc_add_127_23_g191 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_22, A2 => lbl5_en1_count(13), B1 => lbl5_en1_inc_add_127_23_n_22, B2 => lbl5_en1_count(13), ZN => lbl5_en1_n_297);
  lbl5_en1_inc_add_127_23_g192 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_22, B1 => lbl5_en1_count(13), ZN => lbl5_en1_inc_add_127_23_n_24);
  lbl5_en1_inc_add_127_23_g193 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_20, A2 => lbl5_en1_count(12), B1 => lbl5_en1_inc_add_127_23_n_20, B2 => lbl5_en1_count(12), ZN => lbl5_en1_n_296);
  lbl5_en1_inc_add_127_23_g194 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_20, B1 => lbl5_en1_count(12), ZN => lbl5_en1_inc_add_127_23_n_22);
  lbl5_en1_inc_add_127_23_g195 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_18, A2 => lbl5_en1_count(11), B1 => lbl5_en1_inc_add_127_23_n_18, B2 => lbl5_en1_count(11), ZN => FE_PHN170_lbl5_en1_n_295);
  lbl5_en1_inc_add_127_23_g196 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_18, B1 => lbl5_en1_count(11), ZN => lbl5_en1_inc_add_127_23_n_20);
  lbl5_en1_inc_add_127_23_g197 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_16, A2 => lbl5_en1_count(10), B1 => lbl5_en1_inc_add_127_23_n_16, B2 => lbl5_en1_count(10), ZN => lbl5_en1_n_294);
  lbl5_en1_inc_add_127_23_g198 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_16, B1 => lbl5_en1_count(10), ZN => lbl5_en1_inc_add_127_23_n_18);
  lbl5_en1_inc_add_127_23_g199 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_14, A2 => lbl5_en1_count(9), B1 => lbl5_en1_inc_add_127_23_n_14, B2 => lbl5_en1_count(9), ZN => lbl5_en1_n_293);
  lbl5_en1_inc_add_127_23_g200 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_14, B1 => lbl5_en1_count(9), ZN => lbl5_en1_inc_add_127_23_n_16);
  lbl5_en1_inc_add_127_23_g201 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_12, A2 => lbl5_en1_count(8), B1 => lbl5_en1_inc_add_127_23_n_12, B2 => lbl5_en1_count(8), ZN => lbl5_en1_n_292);
  lbl5_en1_inc_add_127_23_g202 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_12, B1 => lbl5_en1_count(8), ZN => lbl5_en1_inc_add_127_23_n_14);
  lbl5_en1_inc_add_127_23_g203 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_10, A2 => lbl5_en1_count(7), B1 => lbl5_en1_inc_add_127_23_n_10, B2 => lbl5_en1_count(7), ZN => lbl5_en1_n_291);
  lbl5_en1_inc_add_127_23_g204 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_10, B1 => lbl5_en1_count(7), ZN => lbl5_en1_inc_add_127_23_n_12);
  lbl5_en1_inc_add_127_23_g205 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_8, A2 => FE_PHN325_lbl5_en1_count_6, B1 => lbl5_en1_inc_add_127_23_n_8, B2 => lbl5_en1_count(6), ZN => lbl5_en1_n_290);
  lbl5_en1_inc_add_127_23_g206 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_8, B1 => lbl5_en1_count(6), ZN => lbl5_en1_inc_add_127_23_n_10);
  lbl5_en1_inc_add_127_23_g207 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_6, A2 => lbl5_en1_count(5), B1 => lbl5_en1_inc_add_127_23_n_6, B2 => lbl5_en1_count(5), ZN => lbl5_en1_n_289);
  lbl5_en1_inc_add_127_23_g208 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_6, B1 => lbl5_en1_count(5), ZN => lbl5_en1_inc_add_127_23_n_8);
  lbl5_en1_inc_add_127_23_g209 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_4, A2 => lbl5_en1_count(4), B1 => lbl5_en1_inc_add_127_23_n_4, B2 => lbl5_en1_count(4), ZN => lbl5_en1_n_288);
  lbl5_en1_inc_add_127_23_g210 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_4, B1 => lbl5_en1_count(4), ZN => lbl5_en1_inc_add_127_23_n_6);
  lbl5_en1_inc_add_127_23_g211 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_2, A2 => lbl5_en1_count(3), B1 => lbl5_en1_inc_add_127_23_n_2, B2 => lbl5_en1_count(3), ZN => lbl5_en1_n_287);
  lbl5_en1_inc_add_127_23_g212 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_2, B1 => lbl5_en1_count(3), ZN => lbl5_en1_inc_add_127_23_n_4);
  lbl5_en1_inc_add_127_23_g213 : MOAI22D0BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_0, A2 => lbl5_en1_count(2), B1 => lbl5_en1_inc_add_127_23_n_0, B2 => lbl5_en1_count(2), ZN => lbl5_en1_n_286);
  lbl5_en1_inc_add_127_23_g214 : IND2D1BWP7T port map(A1 => lbl5_en1_inc_add_127_23_n_0, B1 => lbl5_en1_count(2), ZN => lbl5_en1_inc_add_127_23_n_2);
  lbl5_en1_inc_add_127_23_g215 : CKXOR2D0BWP7T port map(A1 => lbl5_en1_count(0), A2 => lbl5_en1_count(1), Z => FE_PHN190_lbl5_en1_n_285);
  lbl5_en1_inc_add_127_23_g216 : ND2D1BWP7T port map(A1 => lbl5_en1_count(0), A2 => lbl5_en1_count(1), ZN => lbl5_en1_inc_add_127_23_n_0);
  lbl2_pxl_g8183 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_208, A2 => lbl2_pxl_n_191, A3 => lbl2_pxl_n_125, A4 => lbl2_pxl_n_104, ZN => lbl2_pixelator_color(2));
  lbl2_pxl_g8184 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_210, A2 => lbl2_pxl_n_191, A3 => lbl2_pxl_n_177, ZN => lbl2_pixelator_color(0));
  lbl2_pxl_g8185 : ND4D0BWP7T port map(A1 => lbl2_pxl_n_207, A2 => lbl2_pxl_n_184, A3 => lbl2_pxl_n_181, A4 => lbl2_pxl_n_185, ZN => lbl2_pxl_n_210);
  lbl2_pxl_g8186 : AN3D0BWP7T port map(A1 => lbl2_pxl_n_206, A2 => lbl2_pxl_n_195, A3 => lbl2_pxl_n_120, Z => lbl2_pixelator_color(3));
  lbl2_pxl_g8187 : ND4D0BWP7T port map(A1 => lbl2_pxl_n_205, A2 => lbl2_pxl_n_195, A3 => lbl2_pxl_n_167, A4 => lbl2_pxl_n_159, ZN => lbl2_pxl_n_208);
  lbl2_pxl_g8188 : AN4D0BWP7T port map(A1 => lbl2_pxl_n_201, A2 => lbl2_pxl_n_194, A3 => lbl2_pxl_n_197, A4 => lbl2_pxl_n_167, Z => lbl2_pxl_n_207);
  lbl2_pxl_g8189 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_203, A2 => lbl2_pxl_n_175, A3 => lbl2_pxl_n_125, ZN => lbl2_pxl_n_206);
  lbl2_pxl_g8190 : AOI211XD0BWP7T port map(A1 => lbl2_pxl_n_176, A2 => position_0(10), B => lbl2_pxl_n_202, C => lbl2_pxl_n_157, ZN => lbl2_pxl_n_205);
  lbl2_pxl_g8191 : AN4D1BWP7T port map(A1 => lbl2_pxl_n_199, A2 => lbl2_pxl_n_195, A3 => lbl2_pxl_n_198, A4 => lbl2_pxl_n_178, Z => lbl2_pixelator_color(1));
  lbl2_pxl_g8192 : ND4D0BWP7T port map(A1 => lbl2_pxl_n_199, A2 => lbl2_pxl_n_184, A3 => lbl2_pxl_n_179, A4 => lbl2_pxl_n_173, ZN => lbl2_pxl_n_203);
  lbl2_pxl_g8193 : OAI31D0BWP7T port map(A1 => lbl2_pxl_n_124, A2 => lbl2_pxl_n_136, A3 => lbl2_pxl_n_183, B => lbl2_pxl_n_200, ZN => lbl2_pxl_n_202);
  lbl2_pxl_g8194 : OA221D0BWP7T port map(A1 => lbl2_pxl_n_193, A2 => lbl2_pxl_n_163, B1 => lbl2_pxl_n_160, B2 => lbl2_pxl_n_187, C => lbl2_pxl_n_186, Z => lbl2_pxl_n_201);
  lbl2_pxl_g8195 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_196, A2 => lbl2_pxl_n_188, A3 => lbl2_pxl_n_180, A4 => lbl2_pxl_n_177, ZN => lbl2_pxl_n_200);
  lbl2_pxl_g8196 : IINR4D0BWP7T port map(A1 => lbl2_pxl_n_181, A2 => lbl2_pxl_n_2, B1 => lbl2_pxl_n_190, B2 => lbl2_pxl_n_180, ZN => lbl2_pxl_n_198);
  lbl2_pxl_g8197 : OA21D0BWP7T port map(A1 => lbl2_pxl_n_193, A2 => lbl2_pxl_n_155, B => lbl2_pxl_n_194, Z => lbl2_pxl_n_199);
  lbl2_pxl_g8198 : IINR4D0BWP7T port map(A1 => lbl2_pxl_n_158, A2 => lbl2_pxl_n_120, B1 => lbl2_pxl_n_189, B2 => lbl2_pxl_n_104, ZN => lbl2_pxl_n_197);
  lbl2_pxl_g8199 : OAI22D0BWP7T port map(A1 => lbl2_pxl_n_193, A2 => lbl2_pxl_n_164, B1 => lbl2_pxl_n_187, B2 => lbl2_pxl_n_149, ZN => lbl2_pxl_n_196);
  lbl2_pxl_g8200 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_193, B1 => lbl2_pxl_n_113, B2 => lbl2_pxl_n_148, ZN => lbl2_pxl_n_195);
  lbl2_pxl_g8201 : IND4D0BWP7T port map(A1 => lbl2_pxl_n_113, B1 => lbl2_pxl_n_116, B2 => lbl2_pxl_n_148, B3 => lbl2_pxl_n_192, ZN => lbl2_pxl_n_194);
  lbl2_pxl_g8202 : INVD1BWP7T port map(I => lbl2_pxl_n_192, ZN => lbl2_pxl_n_193);
  lbl2_pxl_g8203 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_187, A2 => lbl2_pxl_n_150, A3 => lbl2_pxl_n_131, ZN => lbl2_pxl_n_192);
  lbl2_pxl_g8204 : OAI211D1BWP7T port map(A1 => lbl2_pxl_n_88, A2 => lbl2_pxl_n_174, B => lbl2_pxl_n_158, C => lbl2_pxl_n_159, ZN => lbl2_pxl_n_190);
  lbl2_pxl_g8205 : IND4D0BWP7T port map(A1 => lbl2_pxl_n_175, B1 => lbl2_pxl_n_173, B2 => lbl2_pxl_n_178, B3 => lbl2_pxl_n_2, ZN => lbl2_pxl_n_191);
  lbl2_pxl_g8206 : OAI32D1BWP7T port map(A1 => lbl2_pxl_n_126, A2 => lbl2_pxl_n_123, A3 => lbl2_pxl_n_152, B1 => lbl2_pxl_n_111, B2 => lbl2_pxl_n_183, ZN => lbl2_pxl_n_189);
  lbl2_pxl_g8207 : OAI22D0BWP7T port map(A1 => lbl2_pxl_n_183, A2 => lbl2_pxl_n_107, B1 => lbl2_pxl_n_174, B2 => lbl2_pxl_n_112, ZN => lbl2_pxl_n_188);
  lbl2_pxl_g8208 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_183, B1 => lbl2_pxl_n_151, ZN => lbl2_pxl_n_187);
  lbl2_pxl_g8209 : IND4D0BWP7T port map(A1 => lbl2_pxl_n_124, B1 => lbl2_pxl_n_139, B2 => lbl2_pxl_n_136, B3 => lbl2_pxl_n_182, ZN => lbl2_pxl_n_186);
  lbl2_pxl_g8210 : AOI222D0BWP7T port map(A1 => lbl2_pxl_n_170, A2 => position_1(10), B1 => lbl2_pxl_n_165, B2 => lbl2_pxl_n_143, C1 => lbl2_pxl_n_169, C2 => lbl2_pxl_n_147, ZN => lbl2_pxl_n_185);
  lbl2_pxl_g8211 : INVD1BWP7T port map(I => lbl2_pxl_n_182, ZN => lbl2_pxl_n_183);
  lbl2_pxl_g8212 : OR2D1BWP7T port map(A1 => lbl2_pxl_n_174, A2 => lbl2_pxl_n_118, Z => lbl2_pxl_n_184);
  lbl2_pxl_g8213 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_174, A2 => lbl2_pxl_n_142, ZN => lbl2_pxl_n_182);
  lbl2_pxl_g8214 : AO21D0BWP7T port map(A1 => lbl2_pxl_n_112, A2 => lbl2_pxl_n_88, B => lbl2_pxl_n_174, Z => lbl2_pxl_n_179);
  lbl2_pxl_g8215 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_174, B1 => player_state_1(0), B2 => lbl2_pxl_n_115, ZN => lbl2_pxl_n_181);
  lbl2_pxl_g8216 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_174, A2 => lbl2_pxl_n_114, A3 => player_state_1(0), ZN => lbl2_pxl_n_180);
  lbl2_pxl_g8217 : OAI221D0BWP7T port map(A1 => lbl2_pxl_n_166, A2 => lbl2_pxl_n_127, B1 => lbl2_pxl_n_130, B2 => lbl2_pxl_n_161, C => lbl2_pxl_n_168, ZN => lbl2_pxl_n_176);
  lbl2_pxl_g8218 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_172, A2 => lbl2_pxl_n_119, ZN => lbl2_pxl_n_178);
  lbl2_pxl_g8219 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_171, A2 => lbl2_pxl_n_99, ZN => lbl2_pxl_n_177);
  lbl2_pxl_g8220 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_171, A2 => lbl2_pxl_n_119, A3 => lbl2_pxl_n_97, A4 => lbl2_data_synced(7), ZN => lbl2_pxl_n_175);
  lbl2_pxl_g8222 : IND4D0BWP7T port map(A1 => lbl2_pxl_n_119, B1 => lbl2_pxl_n_97, B2 => lbl2_pxl_n_99, B3 => lbl2_pxl_n_172, ZN => lbl2_pxl_n_174);
  lbl2_pxl_g8223 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_147, B1 => lbl2_pxl_n_121, B2 => lbl2_pxl_n_169, ZN => lbl2_pxl_n_173);
  lbl2_pxl_g8224 : INVD0BWP7T port map(I => lbl2_pxl_n_172, ZN => lbl2_pxl_n_171);
  lbl2_pxl_g8225 : OAI22D0BWP7T port map(A1 => lbl2_pxl_n_166, A2 => lbl2_pxl_n_132, B1 => lbl2_pxl_n_161, B2 => lbl2_pxl_n_138, ZN => lbl2_pxl_n_170);
  lbl2_pxl_g8226 : INR3D0BWP7T port map(A1 => lbl2_pxl_n_169, B1 => lbl2_pxl_n_121, B2 => lbl2_pxl_n_147, ZN => lbl2_pxl_n_172);
  lbl2_pxl_g8227 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_131, A2 => position_1(10), B1 => lbl2_pxl_n_128, B2 => position_0(10), C => lbl2_pxl_n_166, ZN => lbl2_pxl_n_169);
  lbl2_pxl_g8228 : AOI32D1BWP7T port map(A1 => lbl2_pxl_n_165, A2 => lbl2_pxl_n_144, A3 => lbl2_pxl_n_134, B1 => lbl2_pxl_n_156, B2 => lbl2_pxl_n_137, ZN => lbl2_pxl_n_168);
  lbl2_pxl_g8229 : IND4D0BWP7T port map(A1 => lbl2_pxl_n_155, B1 => lbl2_pxl_n_100, B2 => lbl2_pxl_n_132, B3 => lbl2_pxl_n_162, ZN => lbl2_pxl_n_167);
  lbl2_pxl_g8230 : OAI211D1BWP7T port map(A1 => lbl2_pxl_n_8, A2 => lbl2_pxl_n_135, B => lbl2_pxl_n_165, C => lbl2_pxl_n_144, ZN => lbl2_pxl_n_166);
  lbl2_pxl_g8231 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_129, A2 => position_0(10), B1 => lbl2_pxl_n_139, B2 => position_1(10), C => lbl2_pxl_n_161, ZN => lbl2_pxl_n_165);
  lbl2_pxl_g8232 : OA31D1BWP7T port map(A1 => lbl2_data_synced(3), A2 => lbl2_pxl_n_100, A3 => lbl2_pxl_n_155, B => lbl2_pxl_n_127, Z => lbl2_pxl_n_164);
  lbl2_pxl_g8233 : MAOI22D0BWP7T port map(A1 => lbl2_pxl_n_127, A2 => lbl2_pxl_n_140, B1 => lbl2_pxl_n_155, B2 => lbl2_pxl_n_106, ZN => lbl2_pxl_n_163);
  lbl2_pxl_g8234 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_154, A2 => lbl2_pxl_n_150, ZN => lbl2_pxl_n_162);
  lbl2_pxl_g8235 : MAOI22D0BWP7T port map(A1 => lbl2_pxl_n_130, A2 => lbl2_pxl_n_133, B1 => lbl2_pxl_n_150, B2 => lbl2_pxl_n_132, ZN => lbl2_pxl_n_160);
  lbl2_pxl_g8236 : OAI211D1BWP7T port map(A1 => lbl2_pxl_n_8, A2 => lbl2_pxl_n_136, B => lbl2_pxl_n_156, C => lbl2_pxl_n_141, ZN => lbl2_pxl_n_161);
  lbl2_pxl_g8237 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_152, A2 => lbl2_pxl_n_141, ZN => lbl2_pxl_n_157);
  lbl2_pxl_g8238 : IND2D1BWP7T port map(A1 => player_state_1(0), B1 => lbl2_pxl_n_153, ZN => lbl2_pxl_n_159);
  lbl2_pxl_g8239 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_153, A2 => player_state_1(0), ZN => lbl2_pxl_n_158);
  lbl2_pxl_g8240 : ND4D0BWP7T port map(A1 => lbl2_pxl_n_151, A2 => lbl2_pxl_n_122, A3 => lbl2_pxl_n_95, A4 => lbl2_pxl_n_87, ZN => lbl2_pxl_n_154);
  lbl2_pxl_g8241 : INR2XD0BWP7T port map(A1 => lbl2_pxl_n_123, B1 => lbl2_pxl_n_152, ZN => lbl2_pxl_n_156);
  lbl2_pxl_g8242 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_113, B1 => lbl2_pxl_n_117, B2 => lbl2_pxl_n_148, ZN => lbl2_pxl_n_155);
  lbl2_pxl_g8243 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_145, A2 => lbl2_pxl_n_109, ZN => lbl2_pxl_n_153);
  lbl2_pxl_g8244 : OAI211D1BWP7T port map(A1 => lbl2_pxl_n_94, A2 => lbl2_pxl_n_54, B => lbl2_pxl_n_146, C => lbl2_pxl_n_109, ZN => lbl2_pxl_n_152);
  lbl2_pxl_g8245 : OA21D0BWP7T port map(A1 => lbl2_pxl_n_135, A2 => lbl2_pxl_n_133, B => lbl2_pxl_n_130, Z => lbl2_pxl_n_149);
  lbl2_pxl_g8246 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_139, A2 => lbl2_pxl_n_137, A3 => lbl2_pxl_n_124, ZN => lbl2_pxl_n_151);
  lbl2_pxl_g8247 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_133, B1 => lbl2_pxl_n_135, B2 => lbl2_pxl_n_130, ZN => lbl2_pxl_n_150);
  lbl2_pxl_g8248 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_140, A2 => lbl2_pxl_n_128, ZN => lbl2_pxl_n_148);
  lbl2_pxl_g8249 : AN2D1BWP7T port map(A1 => lbl2_pxl_n_140, A2 => position_1(10), Z => lbl2_pxl_n_147);
  lbl2_pxl_g8250 : CKND1BWP7T port map(I => lbl2_pxl_n_145, ZN => lbl2_pxl_n_146);
  lbl2_pxl_g8251 : INVD0BWP7T port map(I => lbl2_pxl_n_144, ZN => lbl2_pxl_n_143);
  lbl2_pxl_g8252 : OAI211D1BWP7T port map(A1 => lbl2_pxl_n_111, A2 => lbl2_pxl_n_107, B => lbl2_pxl_n_122, C => lbl2_pxl_n_105, ZN => lbl2_pxl_n_142);
  lbl2_pxl_g8253 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_125, B1 => lbl2_pxl_n_91, B2 => lbl2_pxl_n_120, ZN => lbl2_pxl_n_145);
  lbl2_pxl_g8254 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_133, A2 => position_1(10), ZN => lbl2_pxl_n_144);
  lbl2_pxl_g8255 : INVD0BWP7T port map(I => lbl2_pxl_n_139, ZN => lbl2_pxl_n_138);
  lbl2_pxl_g8256 : INVD0BWP7T port map(I => lbl2_pxl_n_137, ZN => lbl2_pxl_n_136);
  lbl2_pxl_g8257 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_123, A2 => lbl2_pxl_n_126, ZN => lbl2_pxl_n_141);
  lbl2_pxl_g8258 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_108, A2 => lbl2_pxl_n_1, A3 => lbl2_pxl_n_30, ZN => lbl2_pxl_n_140);
  lbl2_pxl_g8259 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_1, A2 => lbl2_pxl_n_103, A3 => lbl2_pxl_n_6, A4 => lbl2_pxl_n_16, ZN => lbl2_pxl_n_139);
  lbl2_pxl_g8260 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_0, A2 => lbl2_pxl_n_103, A3 => lbl2_pxl_n_6, A4 => lbl2_pxl_n_23, ZN => lbl2_pxl_n_137);
  lbl2_pxl_g8261 : INVD0BWP7T port map(I => lbl2_pxl_n_135, ZN => lbl2_pxl_n_134);
  lbl2_pxl_g8262 : INVD1BWP7T port map(I => lbl2_pxl_n_132, ZN => lbl2_pxl_n_131);
  lbl2_pxl_g8263 : INVD1BWP7T port map(I => lbl2_pxl_n_129, ZN => lbl2_pxl_n_130);
  lbl2_pxl_g8264 : INVD0BWP7T port map(I => lbl2_pxl_n_128, ZN => lbl2_pxl_n_127);
  lbl2_pxl_g8265 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_0, B1 => lbl2_pxl_n_20, B2 => lbl2_pxl_n_110, ZN => lbl2_pxl_n_135);
  lbl2_pxl_g8266 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_1, A2 => lbl2_pxl_n_102, A3 => lbl2_dx(3), A4 => lbl2_pxl_n_29, ZN => lbl2_pxl_n_133);
  lbl2_pxl_g8267 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_1, B1 => lbl2_pxl_n_25, B2 => lbl2_pxl_n_110, ZN => lbl2_pxl_n_132);
  lbl2_pxl_g8268 : NR4D0BWP7T port map(A1 => lbl2_pxl_n_0, A2 => lbl2_pxl_n_102, A3 => lbl2_dx(3), A4 => lbl2_pxl_n_27, ZN => lbl2_pxl_n_129);
  lbl2_pxl_g8269 : NR3D0BWP7T port map(A1 => lbl2_pxl_n_108, A2 => lbl2_pxl_n_0, A3 => lbl2_pxl_n_18, ZN => lbl2_pxl_n_128);
  lbl2_pxl_g8270 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_107, A2 => lbl2_pxl_n_8, ZN => lbl2_pxl_n_126);
  lbl2_pxl_g8271 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_112, A2 => lbl2_pxl_n_8, ZN => lbl2_pxl_n_125);
  lbl2_pxl_g8272 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_111, A2 => lbl2_pxl_n_107, ZN => lbl2_pxl_n_124);
  lbl2_pxl_g8273 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_111, B1 => position_1(10), ZN => lbl2_pxl_n_123);
  lbl2_pxl_g8274 : INR3D0BWP7T port map(A1 => lbl2_pxl_n_88, B1 => lbl2_pxl_n_98, B2 => lbl2_pxl_n_96, ZN => lbl2_pxl_n_122);
  lbl2_pxl_g8275 : AOI211D1BWP7T port map(A1 => lbl2_pxl_n_84, A2 => lbl2_pxl_n_77, B => lbl2_pxl_n_15, C => lbl2_pxl_n_8, ZN => lbl2_pxl_n_121);
  lbl2_pxl_g8276 : OR2D1BWP7T port map(A1 => lbl2_pxl_n_118, A2 => lbl2_pxl_n_8, Z => lbl2_pxl_n_120);
  lbl2_pxl_g8277 : AOI211D1BWP7T port map(A1 => lbl2_pxl_n_79, A2 => lbl2_pxl_n_81, B => lbl2_pxl_n_32, C => FE_DBTN22_position_1_10, ZN => lbl2_pxl_n_119);
  lbl2_pxl_g8278 : INVD1BWP7T port map(I => lbl2_pxl_n_116, ZN => lbl2_pxl_n_117);
  lbl2_pxl_g8279 : INVD0BWP7T port map(I => lbl2_pxl_n_114, ZN => lbl2_pxl_n_115);
  lbl2_pxl_g8280 : IND2D1BWP7T port map(A1 => player_state_0(0), B1 => lbl2_pxl_n_96, ZN => lbl2_pxl_n_118);
  lbl2_pxl_g8281 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_82, A2 => lbl2_pxl_n_83, B => lbl2_pxl_n_32, ZN => lbl2_pxl_n_116);
  lbl2_pxl_g8282 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_96, B1 => lbl2_pxl_n_98, ZN => lbl2_pxl_n_114);
  lbl2_pxl_g8283 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_78, A2 => lbl2_pxl_n_80, B => lbl2_pxl_n_15, ZN => lbl2_pxl_n_113);
  lbl2_pxl_g8284 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_96, A2 => player_state_0(0), ZN => lbl2_pxl_n_112);
  lbl2_pxl_g8285 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_101, A2 => lbl2_pxl_n_42, ZN => lbl2_pxl_n_111);
  lbl2_pxl_g8286 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_100, B1 => lbl2_data_synced(3), ZN => lbl2_pxl_n_106);
  lbl2_pxl_g8287 : OAI211D1BWP7T port map(A1 => lbl2_pxl_n_42, A2 => lbl2_pxl_n_43, B => lbl2_pxl_n_93, C => lbl2_pxl_n_37, ZN => lbl2_pxl_n_105);
  lbl2_pxl_g8288 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_90, A2 => lbl2_dy_vec(2), B => lbl2_dy_vec(3), ZN => lbl2_pxl_n_110);
  lbl2_pxl_g8289 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_98, A2 => position_1(10), ZN => lbl2_pxl_n_109);
  lbl2_pxl_g8290 : OAI21D0BWP7T port map(A1 => lbl2_pxl_n_89, A2 => lbl2_dy_vec(2), B => lbl2_dy_vec(3), ZN => lbl2_pxl_n_108);
  lbl2_pxl_g8291 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_101, A2 => lbl2_pxl_n_43, ZN => lbl2_pxl_n_107);
  lbl2_pxl_g8292 : INR2D1BWP7T port map(A1 => lbl2_pxl_n_88, B1 => lbl2_pxl_n_91, ZN => lbl2_pxl_n_104);
  lbl2_pxl_g8293 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_92, A2 => lbl2_dx(2), ZN => lbl2_pxl_n_103);
  lbl2_pxl_g8294 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_92, A2 => lbl2_pxl_n_3, ZN => lbl2_pxl_n_102);
  lbl2_pxl_g8295 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_37, B1 => lbl2_pxl_n_90, ZN => lbl2_pxl_n_101);
  lbl2_pxl_g8296 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_65, A2 => lbl2_walls(3), B1 => lbl2_pxl_n_67, B2 => lbl2_walls(2), C => lbl2_pxl_n_86, ZN => lbl2_pxl_n_100);
  lbl2_pxl_g8298 : AOI222D0BWP7T port map(A1 => lbl2_pxl_n_56, A2 => lbl2_pxl_n_55, B1 => lbl2_pxl_n_70, B2 => lbl2_jumps_synced(0), C1 => lbl2_pxl_n_68, C2 => lbl2_jumps_synced(2), ZN => lbl2_pxl_n_95);
  lbl2_pxl_g8299 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_69, A2 => lbl2_jumps_synced(5), B1 => lbl2_pxl_n_71, B2 => lbl2_jumps_synced(7), C => lbl2_pxl_n_76, ZN => lbl2_pxl_n_99);
  lbl2_pxl_g8300 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_93, A2 => lbl2_pxl_n_37, ZN => lbl2_pxl_n_94);
  lbl2_pxl_g8301 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_61, A2 => lbl2_pxl_n_5, B1 => lbl2_pxl_n_62, B2 => direction_1(0), C => lbl2_pxl_n_32, ZN => lbl2_pxl_n_98);
  lbl2_pxl_g8302 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_60, A2 => lbl2_walls(4), B1 => lbl2_pxl_n_59, B2 => lbl2_walls(6), C => lbl2_pxl_n_85, ZN => lbl2_pxl_n_97);
  lbl2_pxl_g8303 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_61, A2 => lbl2_pxl_n_10, B1 => lbl2_pxl_n_62, B2 => direction_0(0), C => lbl2_pxl_n_15, ZN => lbl2_pxl_n_96);
  lbl2_pxl_g8304 : INVD0BWP7T port map(I => lbl2_pxl_n_90, ZN => lbl2_pxl_n_89);
  lbl2_pxl_g8305 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_75, A2 => lbl2_pxl_n_38, ZN => lbl2_pxl_n_93);
  lbl2_pxl_g8306 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_69, A2 => lbl2_jumps_synced(1), B1 => lbl2_pxl_n_71, B2 => lbl2_jumps_synced(3), ZN => lbl2_pxl_n_87);
  lbl2_pxl_g8307 : AO22D0BWP7T port map(A1 => lbl2_pxl_n_63, A2 => lbl2_walls(1), B1 => lbl2_walls(0), B2 => lbl2_pxl_n_66, Z => lbl2_pxl_n_86);
  lbl2_pxl_g8308 : AO22D0BWP7T port map(A1 => lbl2_pxl_n_57, A2 => lbl2_walls(5), B1 => lbl2_walls(7), B2 => lbl2_pxl_n_58, Z => lbl2_pxl_n_85);
  lbl2_pxl_g8309 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_37, B1 => lbl2_pxl_n_75, ZN => lbl2_pxl_n_92);
  lbl2_pxl_g8310 : AOI221D0BWP7T port map(A1 => lbl2_pxl_n_50, A2 => lbl2_borders_synced(5), B1 => lbl2_pxl_n_52, B2 => lbl2_borders_synced(6), C => lbl2_pxl_n_73, ZN => lbl2_pxl_n_91);
  lbl2_pxl_g8311 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_74, A2 => lbl2_pxl_n_53, ZN => lbl2_pxl_n_90);
  lbl2_pxl_g8312 : AOI221D1BWP7T port map(A1 => lbl2_pxl_n_50, A2 => lbl2_borders_synced(1), B1 => lbl2_pxl_n_52, B2 => lbl2_borders_synced(2), C => lbl2_pxl_n_72, ZN => lbl2_pxl_n_88);
  lbl2_pxl_g8313 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_59, A2 => lbl2_pxl_n_20, B1 => lbl2_pxl_n_58, B2 => lbl2_pxl_n_26, ZN => lbl2_pxl_n_84);
  lbl2_pxl_g8314 : AOI33D1BWP7T port map(A1 => lbl2_pxl_n_66, A2 => lbl2_pxl_n_5, A3 => direction_1(1), B1 => lbl2_pxl_n_63, B2 => direction_1(0), B3 => direction_1(1), ZN => lbl2_pxl_n_83);
  lbl2_pxl_g8315 : MAOI22D0BWP7T port map(A1 => lbl2_pxl_n_67, A2 => lbl2_pxl_n_25, B1 => lbl2_pxl_n_64, B2 => lbl2_pxl_n_29, ZN => lbl2_pxl_n_82);
  lbl2_pxl_g8316 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_57, A2 => lbl2_pxl_n_17, B1 => lbl2_pxl_n_58, B2 => lbl2_pxl_n_28, ZN => lbl2_pxl_n_81);
  lbl2_pxl_g8317 : MAOI22D0BWP7T port map(A1 => lbl2_pxl_n_63, A2 => lbl2_pxl_n_24, B1 => lbl2_pxl_n_64, B2 => lbl2_pxl_n_27, ZN => lbl2_pxl_n_80);
  lbl2_pxl_g8318 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_60, A2 => lbl2_pxl_n_31, B1 => lbl2_pxl_n_59, B2 => lbl2_pxl_n_25, ZN => lbl2_pxl_n_79);
  lbl2_pxl_g8319 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_67, A2 => lbl2_pxl_n_20, B1 => lbl2_pxl_n_66, B2 => lbl2_pxl_n_19, ZN => lbl2_pxl_n_78);
  lbl2_pxl_g8320 : AOI33D1BWP7T port map(A1 => lbl2_pxl_n_60, A2 => lbl2_pxl_n_10, A3 => direction_0(1), B1 => lbl2_pxl_n_57, B2 => direction_0(0), B3 => direction_0(1), ZN => lbl2_pxl_n_77);
  lbl2_pxl_g8321 : AO22D0BWP7T port map(A1 => lbl2_pxl_n_70, A2 => lbl2_jumps_synced(4), B1 => lbl2_jumps_synced(6), B2 => lbl2_pxl_n_68, Z => lbl2_pxl_n_76);
  lbl2_pxl_g8322 : INVD0BWP7T port map(I => lbl2_pxl_n_74, ZN => lbl2_pxl_n_75);
  lbl2_pxl_g8323 : MAOI222D1BWP7T port map(A => lbl2_pxl_n_46, B => lbl2_pxl_n_35, C => lbl2_pxl_n_34, ZN => lbl2_pxl_n_74);
  lbl2_pxl_g8324 : AO22D0BWP7T port map(A1 => lbl2_pxl_n_49, A2 => lbl2_borders_synced(4), B1 => lbl2_borders_synced(7), B2 => lbl2_pxl_n_51, Z => lbl2_pxl_n_73);
  lbl2_pxl_g8325 : AO22D0BWP7T port map(A1 => lbl2_pxl_n_49, A2 => lbl2_borders_synced(0), B1 => lbl2_borders_synced(3), B2 => lbl2_pxl_n_51, Z => lbl2_pxl_n_72);
  lbl2_pxl_g8326 : INVD0BWP7T port map(I => lbl2_pxl_n_64, ZN => lbl2_pxl_n_65);
  lbl2_pxl_g8327 : AO21D0BWP7T port map(A1 => lbl2_pxl_n_39, A2 => lbl2_dy_vec(1), B => lbl2_pxl_n_51, Z => lbl2_pxl_n_71);
  lbl2_pxl_g8328 : AO21D0BWP7T port map(A1 => lbl2_pxl_n_41, A2 => lbl2_dx(1), B => lbl2_pxl_n_49, Z => lbl2_pxl_n_70);
  lbl2_pxl_g8329 : AO21D0BWP7T port map(A1 => lbl2_pxl_n_40, A2 => lbl2_dy_vec(1), B => lbl2_pxl_n_50, Z => lbl2_pxl_n_69);
  lbl2_pxl_g8330 : AO21D0BWP7T port map(A1 => lbl2_pxl_n_44, A2 => lbl2_dx(1), B => lbl2_pxl_n_52, Z => lbl2_pxl_n_68);
  lbl2_pxl_g8331 : IAO21D0BWP7T port map(A1 => lbl2_dy_vec(3), A2 => lbl2_dy_vec(2), B => lbl2_pxl_n_38, ZN => lbl2_pxl_n_67);
  lbl2_pxl_g8332 : AOI21D0BWP7T port map(A1 => lbl2_dy_vec(3), A2 => lbl2_dy_vec(2), B => lbl2_pxl_n_38, ZN => lbl2_pxl_n_66);
  lbl2_pxl_g8333 : OAI21D0BWP7T port map(A1 => lbl2_dx(3), A2 => lbl2_dx(2), B => lbl2_pxl_n_37, ZN => lbl2_pxl_n_64);
  lbl2_pxl_g8334 : OA21D0BWP7T port map(A1 => lbl2_pxl_n_6, A2 => lbl2_pxl_n_3, B => lbl2_pxl_n_37, Z => lbl2_pxl_n_63);
  lbl2_pxl_g8335 : OAI33D1BWP7T port map(A1 => lbl2_dx(0), A2 => lbl2_pxl_n_6, A3 => lbl2_pxl_n_12, B1 => lbl2_pxl_n_9, B2 => lbl2_dx(3), B3 => lbl2_pxl_n_14, ZN => lbl2_pxl_n_56);
  lbl2_pxl_g8336 : OAI33D1BWP7T port map(A1 => lbl2_dy_vec(0), A2 => lbl2_pxl_n_7, A3 => lbl2_pxl_n_13, B1 => lbl2_pxl_n_11, B2 => lbl2_dy_vec(3), B3 => lbl2_pxl_n_22, ZN => lbl2_pxl_n_55);
  lbl2_pxl_g8337 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_42, A2 => position_1(10), B1 => lbl2_pxl_n_43, B2 => position_0(10), ZN => lbl2_pxl_n_54);
  lbl2_pxl_g8338 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_45, A2 => lbl2_pxl_n_37, ZN => lbl2_pxl_n_62);
  lbl2_pxl_g8339 : OR3XD1BWP7T port map(A1 => lbl2_pxl_n_44, A2 => lbl2_pxl_n_41, A3 => lbl2_pxl_n_38, Z => lbl2_pxl_n_61);
  lbl2_pxl_g8340 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_13, A2 => lbl2_dy_vec(3), B => lbl2_pxl_n_47, ZN => lbl2_pxl_n_60);
  lbl2_pxl_g8341 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_22, A2 => lbl2_pxl_n_7, B => lbl2_pxl_n_47, ZN => lbl2_pxl_n_59);
  lbl2_pxl_g8342 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_14, A2 => lbl2_pxl_n_6, B => lbl2_pxl_n_48, ZN => lbl2_pxl_n_58);
  lbl2_pxl_g8343 : AOI21D0BWP7T port map(A1 => lbl2_pxl_n_12, A2 => lbl2_dx(3), B => lbl2_pxl_n_48, ZN => lbl2_pxl_n_57);
  lbl2_pxl_g8344 : INVD0BWP7T port map(I => lbl2_pxl_n_38, ZN => lbl2_pxl_n_53);
  lbl2_pxl_g8345 : AN2D1BWP7T port map(A1 => lbl2_pxl_n_44, A2 => lbl2_dy_vec(0), Z => lbl2_pxl_n_52);
  lbl2_pxl_g8346 : AN2D1BWP7T port map(A1 => lbl2_pxl_n_39, A2 => lbl2_dx(0), Z => lbl2_pxl_n_51);
  lbl2_pxl_g8347 : AN2D1BWP7T port map(A1 => lbl2_pxl_n_40, A2 => lbl2_pxl_n_9, Z => lbl2_pxl_n_50);
  lbl2_pxl_g8348 : AN2D1BWP7T port map(A1 => lbl2_pxl_n_41, A2 => lbl2_pxl_n_11, Z => lbl2_pxl_n_49);
  lbl2_pxl_g8349 : OAI221D0BWP7T port map(A1 => lbl2_dx(2), A2 => lbl2_dx(0), B1 => lbl2_pxl_n_9, B2 => lbl2_pxl_n_3, C => lbl2_pxl_n_36, ZN => lbl2_pxl_n_46);
  lbl2_pxl_g8350 : NR2D0BWP7T port map(A1 => lbl2_pxl_n_40, A2 => lbl2_pxl_n_39, ZN => lbl2_pxl_n_45);
  lbl2_pxl_g8351 : OA22D0BWP7T port map(A1 => lbl2_pxl_n_13, A2 => lbl2_pxl_n_7, B1 => lbl2_dy_vec(3), B2 => lbl2_pxl_n_22, Z => lbl2_pxl_n_48);
  lbl2_pxl_g8352 : OA22D0BWP7T port map(A1 => lbl2_pxl_n_12, A2 => lbl2_pxl_n_6, B1 => lbl2_dx(3), B2 => lbl2_pxl_n_14, Z => lbl2_pxl_n_47);
  lbl2_pxl_g8353 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_22, A2 => lbl2_pxl_n_7, ZN => lbl2_pxl_n_44);
  lbl2_pxl_g8354 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_21, A2 => player_state_0(0), ZN => lbl2_pxl_n_43);
  lbl2_pxl_g8355 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_33, A2 => player_state_1(0), ZN => lbl2_pxl_n_42);
  lbl2_pxl_g8356 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_13, A2 => lbl2_dy_vec(3), ZN => lbl2_pxl_n_41);
  lbl2_pxl_g8359 : MAOI22D0BWP7T port map(A1 => lbl2_dy_vec(2), A2 => lbl2_dy_vec(0), B1 => lbl2_dy_vec(2), B2 => lbl2_dy_vec(0), ZN => lbl2_pxl_n_36);
  lbl2_pxl_g8360 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_12, A2 => lbl2_pxl_n_14, ZN => lbl2_pxl_n_35);
  lbl2_pxl_g8361 : ND2D1BWP7T port map(A1 => lbl2_pxl_n_13, A2 => lbl2_pxl_n_22, ZN => lbl2_pxl_n_34);
  lbl2_pxl_g8362 : NR2XD0BWP7T port map(A1 => lbl2_pxl_n_12, A2 => lbl2_dx(3), ZN => lbl2_pxl_n_40);
  lbl2_pxl_g8363 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_14, A2 => lbl2_pxl_n_6, ZN => lbl2_pxl_n_39);
  lbl2_pxl_g8364 : AOI22D0BWP7T port map(A1 => lbl2_pxl_n_3, A2 => lbl2_dx(3), B1 => lbl2_pxl_n_6, B2 => lbl2_dx(2), ZN => lbl2_pxl_n_38);
  lbl2_pxl_g8365 : MOAI22D0BWP7T port map(A1 => lbl2_pxl_n_7, A2 => lbl2_dy_vec(2), B1 => lbl2_pxl_n_7, B2 => lbl2_dy_vec(2), ZN => lbl2_pxl_n_37);
  lbl2_pxl_g8367 : INVD0BWP7T port map(I => lbl2_pxl_n_30, ZN => lbl2_pxl_n_31);
  lbl2_pxl_g8368 : CKND1BWP7T port map(I => lbl2_pxl_n_28, ZN => lbl2_pxl_n_29);
  lbl2_pxl_g8369 : CKND1BWP7T port map(I => lbl2_pxl_n_26, ZN => lbl2_pxl_n_27);
  lbl2_pxl_g8370 : INVD0BWP7T port map(I => lbl2_pxl_n_23, ZN => lbl2_pxl_n_24);
  lbl2_pxl_g8371 : IND2D1BWP7T port map(A1 => player_state_1(1), B1 => lbl2_n_189, ZN => lbl2_pxl_n_33);
  lbl2_pxl_g8372 : ND2D1BWP7T port map(A1 => lbl2_n_189, A2 => player_state_1(1), ZN => lbl2_pxl_n_32);
  lbl2_pxl_g8373 : CKND2D1BWP7T port map(A1 => lbl2_pxl_n_5, A2 => direction_1(1), ZN => lbl2_pxl_n_30);
  lbl2_pxl_g8374 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_5, A2 => direction_1(1), ZN => lbl2_pxl_n_28);
  lbl2_pxl_g8375 : NR2D1BWP7T port map(A1 => lbl2_pxl_n_10, A2 => direction_0(1), ZN => lbl2_pxl_n_26);
  lbl2_pxl_g8376 : NR2D0BWP7T port map(A1 => direction_1(1), A2 => direction_1(0), ZN => lbl2_pxl_n_25);
  lbl2_pxl_g8377 : CKND2D1BWP7T port map(A1 => direction_0(1), A2 => direction_0(0), ZN => lbl2_pxl_n_23);
  lbl2_pxl_g8378 : ND2D1BWP7T port map(A1 => lbl2_dy_vec(2), A2 => lbl2_dy_vec(1), ZN => lbl2_pxl_n_22);
  lbl2_pxl_g8380 : INVD0BWP7T port map(I => lbl2_pxl_n_18, ZN => lbl2_pxl_n_19);
  lbl2_pxl_g8381 : INVD0BWP7T port map(I => lbl2_pxl_n_16, ZN => lbl2_pxl_n_17);
  lbl2_pxl_g8382 : IND2D1BWP7T port map(A1 => player_state_0(1), B1 => lbl2_n_190, ZN => lbl2_pxl_n_21);
  lbl2_pxl_g8383 : NR2D0BWP7T port map(A1 => direction_0(1), A2 => direction_0(0), ZN => lbl2_pxl_n_20);
  lbl2_pxl_g8384 : CKND2D1BWP7T port map(A1 => lbl2_pxl_n_10, A2 => direction_0(1), ZN => lbl2_pxl_n_18);
  lbl2_pxl_g8385 : CKND2D1BWP7T port map(A1 => direction_1(1), A2 => direction_1(0), ZN => lbl2_pxl_n_16);
  lbl2_pxl_g8386 : ND2D1BWP7T port map(A1 => lbl2_n_190, A2 => player_state_0(1), ZN => lbl2_pxl_n_15);
  lbl2_pxl_g8387 : ND2D1BWP7T port map(A1 => lbl2_dx(1), A2 => lbl2_dx(2), ZN => lbl2_pxl_n_14);
  lbl2_pxl_g8388 : OR2D1BWP7T port map(A1 => lbl2_dy_vec(1), A2 => lbl2_dy_vec(2), Z => lbl2_pxl_n_13);
  lbl2_pxl_g8389 : OR2D1BWP7T port map(A1 => lbl2_dx(1), A2 => lbl2_dx(2), Z => lbl2_pxl_n_12);
  lbl2_pxl_g8390 : INVD1BWP7T port map(I => lbl2_dy_vec(0), ZN => lbl2_pxl_n_11);
  lbl2_pxl_g8391 : INVD1BWP7T port map(I => direction_0(0), ZN => lbl2_pxl_n_10);
  lbl2_pxl_g8392 : INVD0BWP7T port map(I => lbl2_dx(0), ZN => lbl2_pxl_n_9);
  lbl2_pxl_g8393 : INVD1BWP7T port map(I => position_0(10), ZN => lbl2_pxl_n_8);
  lbl2_pxl_g8394 : INVD1BWP7T port map(I => lbl2_dy_vec(3), ZN => lbl2_pxl_n_7);
  lbl2_pxl_g8395 : INVD1BWP7T port map(I => lbl2_dx(3), ZN => lbl2_pxl_n_6);
  lbl2_pxl_g8396 : INVD1BWP7T port map(I => direction_1(0), ZN => lbl2_pxl_n_5);
  lbl2_pxl_g8398 : INVD1BWP7T port map(I => lbl2_dx(2), ZN => lbl2_pxl_n_3);
  lbl2_pxl_g2 : IND3D1BWP7T port map(A1 => lbl2_pxl_n_97, B1 => lbl2_pxl_n_172, B2 => lbl2_data_synced(7), ZN => lbl2_pxl_n_2);
  lbl2_pxl_g8399 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_33, B1 => player_state_1(0), ZN => lbl2_pxl_n_1);
  lbl2_pxl_g8400 : IND2D1BWP7T port map(A1 => lbl2_pxl_n_21, B1 => player_state_0(0), ZN => lbl2_pxl_n_0);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1075 : AN4D1BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_34, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_31, A3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_30, A4 => lbl5_en1_csa_tree_lt_140_15_groupi_n_28, Z => lbl5_en1_n_284);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1076 : AOI31D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_27, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_37, A3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_54, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_33, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_34);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1077 : ND4D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_32, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_24, A3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_21, A4 => lbl5_en1_csa_tree_lt_140_15_groupi_n_23, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_33);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1078 : IND3D0BWP7T port map(A1 => lbl5_en1_n_305, B1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_36, B2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_29, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_32);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1079 : OAI211D1BWP7T port map(A1 => FE_DBTN8_lbl5_en1_n_305, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_36, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_29, C => lbl5_en1_csa_tree_lt_140_15_groupi_n_4, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_31);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1080 : AOI33D1BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_26, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_38, A3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_55, B1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_20, B2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_41, B3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_58, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_30);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1081 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_37, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_54, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_27, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_29);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1082 : AOI33D1BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_25, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_39, A3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_56, B1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_22, B2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_40, B3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_57, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_28);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1083 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_38, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_55, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_26, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_27);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1084 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_39, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_56, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_25, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_26);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1085 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_40, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_57, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_22, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_25);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1086 : AOI33D1BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_18, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_42, A3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_59, B1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_13, B2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_45, B3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_62, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_24);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1087 : AOI31D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_8, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_49, A3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_66, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_19, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_23);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1088 : AOI33D1BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_16, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_43, A3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_60, B1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_12, B2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_46, B3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_63, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_21);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1089 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_41, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_58, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_20, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_22);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1090 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_42, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_59, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_18, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_20);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1091 : ND4D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_17, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_14, A3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_10, A4 => lbl5_en1_csa_tree_lt_140_15_groupi_n_6, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_19);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1092 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_43, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_60, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_16, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_18);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1093 : ND3D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_15, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_44, A3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_61, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_17);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1094 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_44, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_61, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_15, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_16);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1095 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_45, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_62, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_13, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_15);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1096 : AOI33D1BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_11, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_47, A3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_64, B1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_9, B2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_48, B3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_65, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_14);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1097 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_46, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_63, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_12, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_13);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1098 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_47, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_64, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_11, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_12);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1099 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_48, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_65, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_9, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_11);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1100 : AOI33D1BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_7, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_50, A3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_67, B1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_5, B2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_51, B3 => lbl5_en1_csa_tree_lt_140_15_groupi_n_68, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_10);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1101 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_49, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_66, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_8, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_9);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1102 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_50, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_67, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_7, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_8);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1103 : OA21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_51, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_68, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_5, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_7);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1104 : AOI22D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_3, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_52, B1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_53, B2 => lbl5_en1_count(18), ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_6);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1105 : AO21D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_2, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_52, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_3, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_5);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1106 : MAOI222D1BWP7T port map(A => lbl5_en1_n_304, B => lbl5_en1_n_303, C => lbl5_en1_csa_tree_lt_140_15_groupi_n_0, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_4);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1107 : AN2D0BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_2, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_69, Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_3);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1108 : OR2D1BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_53, A2 => lbl5_en1_count(18), Z => lbl5_en1_csa_tree_lt_140_15_groupi_n_2);
  lbl5_en1_csa_tree_lt_140_15_groupi_g1110 : CKND1BWP7T port map(I => lbl5_en1_count(0), ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_0);
  lbl5_en1_csa_tree_lt_140_15_groupi_g882 : FA1D0BWP7T port map(A => lbl5_en1_csa_tree_lt_140_15_groupi_n_124, B => lbl5_en1_count(16), CI => lbl5_en1_csa_tree_lt_140_15_groupi_n_112, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_69, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_51);
  lbl5_en1_csa_tree_lt_140_15_groupi_g883 : FA1D0BWP7T port map(A => lbl5_en1_csa_tree_lt_140_15_groupi_n_112, B => lbl5_en1_count(15), CI => lbl5_en1_csa_tree_lt_140_15_groupi_n_123, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_68, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_50);
  lbl5_en1_csa_tree_lt_140_15_groupi_g884 : FA1D0BWP7T port map(A => lbl5_en1_csa_tree_lt_140_15_groupi_n_121, B => lbl5_en1_count(13), CI => lbl5_en1_csa_tree_lt_140_15_groupi_n_119, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_66, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_48);
  lbl5_en1_csa_tree_lt_140_15_groupi_g885 : FA1D0BWP7T port map(A => FE_DBTN0_lbl5_en1_n_306, B => lbl5_en1_count(2), CI => FE_DBTN8_lbl5_en1_n_305, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_55, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_37);
  lbl5_en1_csa_tree_lt_140_15_groupi_g886 : FA1D0BWP7T port map(A => FE_DBTN3_lbl5_en1_n_307, B => lbl5_en1_count(3), CI => FE_DBTN0_lbl5_en1_n_306, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_56, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_38);
  lbl5_en1_csa_tree_lt_140_15_groupi_g887 : FA1D0BWP7T port map(A => FE_DBTN7_lbl5_en1_n_308, B => lbl5_en1_count(4), CI => FE_DBTN3_lbl5_en1_n_307, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_57, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_39);
  lbl5_en1_csa_tree_lt_140_15_groupi_g888 : FA1D0BWP7T port map(A => FE_DBTN5_lbl5_en1_n_309, B => lbl5_en1_count(5), CI => FE_DBTN7_lbl5_en1_n_308, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_58, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_40);
  lbl5_en1_csa_tree_lt_140_15_groupi_g889 : FA1D0BWP7T port map(A => FE_DBTN6_lbl5_en1_n_310, B => lbl5_en1_count(6), CI => FE_DBTN5_lbl5_en1_n_309, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_59, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_41);
  lbl5_en1_csa_tree_lt_140_15_groupi_g890 : FA1D0BWP7T port map(A => lbl5_en1_csa_tree_lt_140_15_groupi_n_118, B => lbl5_en1_count(7), CI => FE_DBTN6_lbl5_en1_n_310, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_60, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_42);
  lbl5_en1_csa_tree_lt_140_15_groupi_g891 : FA1D0BWP7T port map(A => FE_DBTN4_lbl5_en1_n_313, B => lbl5_en1_count(9), CI => FE_DBTN2_lbl5_en1_n_312, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_62, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_44);
  lbl5_en1_csa_tree_lt_140_15_groupi_g892 : FA1D0BWP7T port map(A => FE_DBTN2_lbl5_en1_n_312, B => lbl5_en1_count(8), CI => lbl5_en1_csa_tree_lt_140_15_groupi_n_118, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_61, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_43);
  lbl5_en1_csa_tree_lt_140_15_groupi_g893 : FA1D0BWP7T port map(A => lbl5_en1_csa_tree_lt_140_15_groupi_n_120, B => lbl5_en1_count(10), CI => FE_DBTN4_lbl5_en1_n_313, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_63, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_45);
  lbl5_en1_csa_tree_lt_140_15_groupi_g894 : FA1D0BWP7T port map(A => FE_DBTN1_lbl5_en1_n_315, B => lbl5_en1_count(11), CI => lbl5_en1_csa_tree_lt_140_15_groupi_n_120, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_64, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_46);
  lbl5_en1_csa_tree_lt_140_15_groupi_g895 : FA1D0BWP7T port map(A => lbl5_en1_csa_tree_lt_140_15_groupi_n_119, B => lbl5_en1_count(12), CI => FE_DBTN1_lbl5_en1_n_315, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_65, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_47);
  lbl5_en1_csa_tree_lt_140_15_groupi_g896 : FA1D0BWP7T port map(A => lbl5_en1_csa_tree_lt_140_15_groupi_n_123, B => lbl5_en1_count(14), CI => lbl5_en1_csa_tree_lt_140_15_groupi_n_121, CO => lbl5_en1_csa_tree_lt_140_15_groupi_n_67, S => lbl5_en1_csa_tree_lt_140_15_groupi_n_49);
  lbl5_en1_csa_tree_lt_140_15_groupi_g897 : OAI21D0BWP7T port map(A1 => lbl5_en1_n_304, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_114, B => lbl5_en1_csa_tree_lt_140_15_groupi_n_54, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_36);
  lbl5_en1_csa_tree_lt_140_15_groupi_g898 : IOA21D1BWP7T port map(A1 => lbl5_en1_csa_tree_lt_140_15_groupi_n_124, A2 => lbl5_en1_count(17), B => lbl5_en1_csa_tree_lt_140_15_groupi_n_53, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_52);
  lbl5_en1_csa_tree_lt_140_15_groupi_g899 : ND2D1BWP7T port map(A1 => lbl5_en1_n_304, A2 => lbl5_en1_csa_tree_lt_140_15_groupi_n_114, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_54);
  lbl5_en1_csa_tree_lt_140_15_groupi_g900 : IND2D1BWP7T port map(A1 => lbl5_en1_count(17), B1 => lbl5_en1_n_320, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_53);
  lbl5_en1_csa_tree_lt_140_15_groupi_g901 : INVD1BWP7T port map(I => lbl5_en1_n_320, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_124);
  lbl5_en1_csa_tree_lt_140_15_groupi_g902 : INVD0BWP7T port map(I => lbl5_en1_n_318, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_123);
  lbl5_en1_csa_tree_lt_140_15_groupi_g904 : INVD1BWP7T port map(I => lbl5_en1_n_317, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_121);
  lbl5_en1_csa_tree_lt_140_15_groupi_g905 : INVD1BWP7T port map(I => lbl5_en1_n_314, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_120);
  lbl5_en1_csa_tree_lt_140_15_groupi_g906 : INVD1BWP7T port map(I => lbl5_en1_n_316, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_119);
  lbl5_en1_csa_tree_lt_140_15_groupi_g907 : INVD1BWP7T port map(I => lbl5_en1_n_311, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_118);
  lbl5_en1_csa_tree_lt_140_15_groupi_g911 : CKND1BWP7T port map(I => lbl5_en1_count(1), ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_114);
  lbl5_en1_csa_tree_lt_140_15_groupi_g913 : INVD1BWP7T port map(I => lbl5_en1_n_319, ZN => lbl5_en1_csa_tree_lt_140_15_groupi_n_112);
  lbl2_sdb_g8558 : OR2D1BWP7T port map(A1 => lbl2_sidebar_color(1), A2 => lbl2_sdb_n_173, Z => lbl2_sidebar_color(0));
  lbl2_sdb_g8559 : OR2D1BWP7T port map(A1 => lbl2_sidebar_color(3), A2 => lbl2_sdb_n_173, Z => lbl2_sidebar_color(2));
  lbl2_sdb_g8560 : INR2D1BWP7T port map(A1 => lbl2_h_count(9), B1 => lbl2_sdb_n_194, ZN => lbl2_sidebar_color(3));
  lbl2_sdb_g8561 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_194, A2 => lbl2_h_count(9), ZN => lbl2_sidebar_color(1));
  lbl2_sdb_g8562 : AOI31D0BWP7T port map(A1 => lbl2_sdb_n_184, A2 => game_state(2), A3 => game_state(0), B => lbl2_sdb_n_193, ZN => lbl2_sdb_n_194);
  lbl2_sdb_g8563 : AO211D0BWP7T port map(A1 => lbl2_sdb_n_168, A2 => lbl2_n_151, B => lbl2_sdb_n_192, C => lbl2_sdb_n_190, Z => lbl2_sdb_n_193);
  lbl2_sdb_g8564 : OAI31D0BWP7T port map(A1 => lbl2_v_count(7), A2 => lbl2_v_count(8), A3 => lbl2_sdb_n_191, B => lbl2_sdb_n_188, ZN => lbl2_sdb_n_192);
  lbl2_sdb_g8565 : OAI21D0BWP7T port map(A1 => lbl2_sdb_n_189, A2 => lbl2_sdb_n_178, B => lbl2_sdb_n_13, ZN => lbl2_sdb_n_191);
  lbl2_sdb_g8566 : OAI31D0BWP7T port map(A1 => lbl2_v_count(7), A2 => lbl2_sdb_n_46, A3 => lbl2_sdb_n_186, B => lbl2_sdb_n_181, ZN => lbl2_sdb_n_190);
  lbl2_sdb_g8567 : OAI32D1BWP7T port map(A1 => lbl2_sdb_n_214, A2 => lbl2_sdb_n_63, A3 => lbl2_sdb_n_169, B1 => lbl2_sdb_n_100, B2 => lbl2_sdb_n_187, ZN => lbl2_sdb_n_189);
  lbl2_sdb_g8568 : IND3D1BWP7T port map(A1 => lbl2_sdb_n_185, B1 => lbl2_v_count(6), B2 => lbl2_v_count(8), ZN => lbl2_sdb_n_188);
  lbl2_sdb_g8569 : OAI222D0BWP7T port map(A1 => lbl2_sdb_n_182, A2 => lbl2_sdb_n_157, B1 => lbl2_sdb_n_10, B2 => lbl2_sdb_n_0, C1 => lbl2_h_count(9), C2 => lbl2_sdb_n_41, ZN => lbl2_sdb_n_187);
  lbl2_sdb_g8570 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_183, A2 => lbl2_sdb_n_31, ZN => lbl2_sdb_n_186);
  lbl2_sdb_g8571 : IND4D0BWP7T port map(A1 => lbl2_sdb_n_100, B1 => lbl2_sdb_n_46, B2 => lbl2_sdb_n_31, B3 => lbl2_sdb_n_180, ZN => lbl2_sdb_n_185);
  lbl2_sdb_g8572 : AN4D0BWP7T port map(A1 => lbl2_sdb_n_174, A2 => lbl2_sdb_n_32, A3 => lbl2_sdb_n_48, A4 => lbl2_n_154, Z => lbl2_sdb_n_184);
  lbl2_sdb_g8573 : OAI22D0BWP7T port map(A1 => lbl2_sdb_n_179, A2 => lbl2_h_count(9), B1 => lbl2_sdb_n_160, B2 => lbl2_sdb_n_10, ZN => lbl2_sdb_n_183);
  lbl2_sdb_g8574 : OAI211D1BWP7T port map(A1 => lbl2_sdb_n_35, A2 => lbl2_sdb_n_107, B => lbl2_sdb_n_177, C => lbl2_sdb_n_141, ZN => lbl2_sdb_n_182);
  lbl2_sdb_g8575 : IOA21D0BWP7T port map(A1 => lbl2_sdb_n_172, A2 => lbl2_sdb_n_143, B => lbl2_sdb_n_176, ZN => lbl2_sdb_n_181);
  lbl2_sdb_g8576 : OAI31D0BWP7T port map(A1 => lbl2_sdb_n_27, A2 => lbl2_sdb_n_107, A3 => lbl2_sdb_n_121, B => lbl2_sdb_n_175, ZN => lbl2_sdb_n_180);
  lbl2_sdb_g8577 : AOI32D1BWP7T port map(A1 => lbl2_sdb_n_155, A2 => lbl2_sdb_n_99, A3 => lbl2_sdb_n_27, B1 => lbl2_sdb_n_171, B2 => lbl2_sdb_n_57, ZN => lbl2_sdb_n_179);
  lbl2_sdb_g8578 : NR4D0BWP7T port map(A1 => lbl2_sdb_n_164, A2 => lbl2_sdb_n_100, A3 => lbl2_sdb_n_16, A4 => game_state(1), ZN => lbl2_sdb_n_178);
  lbl2_sdb_g8579 : AOI222D0BWP7T port map(A1 => lbl2_sdb_n_165, A2 => lbl2_sdb_n_27, B1 => lbl2_sdb_n_125, B2 => lbl2_sdb_n_70, C1 => lbl2_sdb_n_153, C2 => lbl2_sdb_n_12, ZN => lbl2_sdb_n_177);
  lbl2_sdb_g8580 : OAI31D0BWP7T port map(A1 => lbl2_sdb_n_8, A2 => lbl2_sdb_n_2, A3 => lbl2_sdb_n_67, B => lbl2_sdb_n_172, ZN => lbl2_sdb_n_176);
  lbl2_sdb_g8581 : MAOI22D0BWP7T port map(A1 => lbl2_sdb_n_167, A2 => lbl2_sdb_n_72, B1 => lbl2_sdb_n_154, B2 => lbl2_sdb_n_103, ZN => lbl2_sdb_n_175);
  lbl2_sdb_g8582 : OAI211D1BWP7T port map(A1 => lbl2_sdb_n_106, A2 => lbl2_sdb_n_90, B => lbl2_sdb_n_170, C => lbl2_sdb_n_95, ZN => lbl2_sdb_n_174);
  lbl2_sdb_g8583 : INR2D1BWP7T port map(A1 => lbl2_sdb_n_168, B1 => lbl2_n_151, ZN => lbl2_sdb_n_173);
  lbl2_sdb_g8584 : AOI31D0BWP7T port map(A1 => lbl2_sdb_n_158, A2 => lbl2_sdb_n_150, A3 => lbl2_sdb_n_135, B => lbl2_sdb_n_100, ZN => lbl2_sdb_n_171);
  lbl2_sdb_g8585 : ND4D0BWP7T port map(A1 => lbl2_sdb_n_162, A2 => lbl2_sdb_n_24, A3 => lbl2_v_count(8), A4 => lbl2_v_count(7), ZN => lbl2_sdb_n_172);
  lbl2_sdb_g8586 : AOI31D0BWP7T port map(A1 => lbl2_sdb_n_53, A2 => lbl2_sdb_n_19, A3 => lbl2_sdb_n_93, B => lbl2_sdb_n_163, ZN => lbl2_sdb_n_170);
  lbl2_sdb_g8587 : AOI211XD0BWP7T port map(A1 => lbl2_sdb_n_129, A2 => lbl2_sdb_n_14, B => lbl2_sdb_n_166, C => lbl2_sdb_n_124, ZN => lbl2_sdb_n_169);
  lbl2_sdb_g8588 : AOI22D0BWP7T port map(A1 => lbl2_sdb_n_159, A2 => lbl2_sdb_n_109, B1 => lbl2_sdb_n_136, B2 => lbl2_sdb_n_57, ZN => lbl2_sdb_n_167);
  lbl2_sdb_g8589 : AOI211D1BWP7T port map(A1 => lbl2_sdb_n_148, A2 => lbl2_sdb_n_104, B => lbl2_sdb_n_32, C => lbl2_sdb_n_47, ZN => lbl2_sdb_n_168);
  lbl2_sdb_g8590 : OAI221D0BWP7T port map(A1 => lbl2_sdb_n_130, A2 => lbl2_h_count(2), B1 => lbl2_sdb_n_78, B2 => lbl2_sdb_n_115, C => lbl2_sdb_n_161, ZN => lbl2_sdb_n_166);
  lbl2_sdb_g8591 : OAI211D1BWP7T port map(A1 => lbl2_sdb_n_87, A2 => lbl2_sdb_n_121, B => lbl2_sdb_n_150, C => lbl2_sdb_n_136, ZN => lbl2_sdb_n_165);
  lbl2_sdb_g8592 : NR2XD0BWP7T port map(A1 => lbl2_sdb_n_156, A2 => lbl2_sdb_n_146, ZN => lbl2_sdb_n_164);
  lbl2_sdb_g8593 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_149, A2 => lbl2_sdb_n_131, B => lbl2_sdb_n_57, ZN => lbl2_sdb_n_163);
  lbl2_sdb_g8594 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_138, A2 => lbl2_sdb_n_91, B => lbl2_sdb_n_18, ZN => lbl2_sdb_n_162);
  lbl2_sdb_g8595 : OAI21D0BWP7T port map(A1 => lbl2_sdb_n_140, A2 => lbl2_sdb_n_129, B => lbl2_h_count(2), ZN => lbl2_sdb_n_161);
  lbl2_sdb_g8596 : AOI221D0BWP7T port map(A1 => lbl2_sdb_n_92, A2 => lbl2_sdb_n_93, B1 => lbl2_sdb_n_38, B2 => lbl2_sdb_n_70, C => lbl2_sdb_n_152, ZN => lbl2_sdb_n_160);
  lbl2_sdb_g8597 : OA211D0BWP7T port map(A1 => lbl2_sdb_n_23, A2 => lbl2_sdb_n_107, B => lbl2_sdb_n_147, C => lbl2_sdb_n_137, Z => lbl2_sdb_n_159);
  lbl2_sdb_g8598 : AOI31D0BWP7T port map(A1 => lbl2_sdb_n_98, A2 => lbl2_sdb_n_87, A3 => lbl2_sdb_n_54, B => lbl2_sdb_n_145, ZN => lbl2_sdb_n_158);
  lbl2_sdb_g8599 : AOI211D1BWP7T port map(A1 => lbl2_sdb_n_134, A2 => lbl2_sdb_n_117, B => lbl2_sdb_n_27, C => lbl2_v_count(2), ZN => lbl2_sdb_n_157);
  lbl2_sdb_g8600 : OAI31D0BWP7T port map(A1 => lbl2_sdb_n_77, A2 => lbl2_sdb_n_87, A3 => lbl2_sdb_n_119, B => lbl2_sdb_n_151, ZN => lbl2_sdb_n_156);
  lbl2_sdb_g8601 : OAI22D0BWP7T port map(A1 => lbl2_sdb_n_133, A2 => lbl2_sdb_n_116, B1 => lbl2_sdb_n_134, B2 => lbl2_v_count(2), ZN => lbl2_sdb_n_155);
  lbl2_sdb_g8602 : AOI221D0BWP7T port map(A1 => lbl2_sdb_n_118, A2 => lbl2_sdb_n_57, B1 => lbl2_sdb_n_98, B2 => lbl2_sdb_n_28, C => lbl2_sdb_n_120, ZN => lbl2_sdb_n_154);
  lbl2_sdb_g8603 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_144, A2 => lbl2_sdb_n_108, ZN => lbl2_sdb_n_153);
  lbl2_sdb_g8604 : OAI21D0BWP7T port map(A1 => lbl2_sdb_n_29, A2 => lbl2_sdb_n_106, B => lbl2_sdb_n_139, ZN => lbl2_sdb_n_152);
  lbl2_sdb_g8605 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_127, A2 => lbl2_sdb_n_118, B => lbl2_sdb_n_126, ZN => lbl2_sdb_n_151);
  lbl2_sdb_g8606 : AOI222D0BWP7T port map(A1 => lbl2_sdb_n_112, A2 => lbl2_sdb_n_37, B1 => lbl2_sdb_n_82, B2 => lbl2_sdb_n_20, C1 => lbl2_sdb_n_55, C2 => lbl2_sdb_n_93, ZN => lbl2_sdb_n_149);
  lbl2_sdb_g8607 : OA222D0BWP7T port map(A1 => lbl2_sdb_n_113, A2 => lbl2_sdb_n_57, B1 => lbl2_sdb_n_106, B2 => lbl2_sdb_n_80, C1 => lbl2_sdb_n_108, C2 => lbl2_sdb_n_36, Z => lbl2_sdb_n_148);
  lbl2_sdb_g8608 : AOI31D0BWP7T port map(A1 => lbl2_sdb_n_122, A2 => lbl2_sdb_n_102, A3 => lbl2_v_count(2), B => lbl2_sdb_n_142, ZN => lbl2_sdb_n_147);
  lbl2_sdb_g8609 : OAI22D0BWP7T port map(A1 => lbl2_sdb_n_132, A2 => lbl2_sdb_n_106, B1 => lbl2_sdb_n_135, B2 => lbl2_sdb_n_73, ZN => lbl2_sdb_n_146);
  lbl2_sdb_g8610 : OAI22D0BWP7T port map(A1 => lbl2_sdb_n_132, A2 => lbl2_sdb_n_93, B1 => lbl2_sdb_n_114, B2 => lbl2_sdb_n_98, ZN => lbl2_sdb_n_145);
  lbl2_sdb_g8611 : AOI33D1BWP7T port map(A1 => lbl2_sdb_n_118, A2 => lbl2_sdb_n_86, A3 => lbl2_v_count(2), B1 => lbl2_sdb_n_77, B2 => lbl2_sdb_n_14, B3 => lbl2_sdb_n_8, ZN => lbl2_sdb_n_150);
  lbl2_sdb_g8612 : AOI31D0BWP7T port map(A1 => lbl2_sdb_n_97, A2 => lbl2_sdb_n_87, A3 => lbl2_sdb_n_34, B => lbl2_sdb_n_122, ZN => lbl2_sdb_n_144);
  lbl2_sdb_g8613 : AOI31D0BWP7T port map(A1 => lbl2_sdb_n_1, A2 => lbl2_sdb_n_71, A3 => lbl2_n_152, B => lbl2_sdb_n_128, ZN => lbl2_sdb_n_143);
  lbl2_sdb_g8614 : NR2D0BWP7T port map(A1 => lbl2_sdb_n_133, A2 => lbl2_sdb_n_86, ZN => lbl2_sdb_n_142);
  lbl2_sdb_g8615 : IND4D0BWP7T port map(A1 => lbl2_sdb_n_102, B1 => lbl2_v_count(2), B2 => lbl2_sdb_n_70, B3 => lbl2_sdb_n_98, ZN => lbl2_sdb_n_141);
  lbl2_sdb_g8616 : AO33D0BWP7T port map(A1 => lbl2_sdb_n_88, A2 => lbl2_sdb_n_94, A3 => lbl2_sdb_n_8, B1 => lbl2_sdb_n_89, B2 => lbl2_sdb_n_78, B3 => lbl2_sdb_n_12, Z => lbl2_sdb_n_140);
  lbl2_sdb_g8617 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_65, A2 => lbl2_sdb_n_110, B => lbl2_sdb_n_123, ZN => lbl2_sdb_n_139);
  lbl2_sdb_g8618 : OAI21D0BWP7T port map(A1 => lbl2_sdb_n_17, A2 => lbl2_sdb_n_13, B => lbl2_sdb_n_128, ZN => lbl2_sdb_n_138);
  lbl2_sdb_g8619 : MOAI22D0BWP7T port map(A1 => lbl2_sdb_n_120, A2 => lbl2_sdb_n_93, B1 => lbl2_sdb_n_121, B2 => lbl2_sdb_n_93, ZN => lbl2_sdb_n_137);
  lbl2_sdb_g8620 : OAI22D0BWP7T port map(A1 => lbl2_sdb_n_105, A2 => lbl2_sdb_n_25, B1 => lbl2_sdb_n_37, B2 => lbl2_sdb_n_19, ZN => lbl2_sdb_n_131);
  lbl2_sdb_g8621 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_111, A2 => lbl2_sdb_n_88, ZN => lbl2_sdb_n_130);
  lbl2_sdb_g8622 : IND2D1BWP7T port map(A1 => lbl2_sdb_n_107, B1 => lbl2_sdb_n_118, ZN => lbl2_sdb_n_136);
  lbl2_sdb_g8623 : IND2D1BWP7T port map(A1 => lbl2_sdb_n_102, B1 => lbl2_sdb_n_122, ZN => lbl2_sdb_n_135);
  lbl2_sdb_g8624 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_122, A2 => lbl2_sdb_n_77, ZN => lbl2_sdb_n_134);
  lbl2_sdb_g8625 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_118, A2 => lbl2_sdb_n_14, ZN => lbl2_sdb_n_133);
  lbl2_sdb_g8626 : NR2XD0BWP7T port map(A1 => lbl2_sdb_n_120, A2 => lbl2_sdb_n_118, ZN => lbl2_sdb_n_132);
  lbl2_sdb_g8627 : OAI22D0BWP7T port map(A1 => lbl2_sdb_n_109, A2 => lbl2_sdb_n_57, B1 => lbl2_sdb_n_77, B2 => lbl2_sdb_n_11, ZN => lbl2_sdb_n_127);
  lbl2_sdb_g8628 : IAO21D0BWP7T port map(A1 => lbl2_sdb_n_101, A2 => lbl2_sdb_n_110, B => lbl2_sdb_n_121, ZN => lbl2_sdb_n_126);
  lbl2_sdb_g8629 : OAI21D0BWP7T port map(A1 => lbl2_sdb_n_98, A2 => lbl2_sdb_n_87, B => lbl2_sdb_n_103, ZN => lbl2_sdb_n_125);
  lbl2_sdb_g8630 : NR4D0BWP7T port map(A1 => lbl2_sdb_n_89, A2 => lbl2_sdb_n_78, A3 => lbl2_sdb_n_60, A4 => lbl2_sdb_n_11, ZN => lbl2_sdb_n_124);
  lbl2_sdb_g8631 : OAI22D0BWP7T port map(A1 => lbl2_sdb_n_74, A2 => lbl2_sdb_n_108, B1 => lbl2_sdb_n_85, B2 => lbl2_sdb_n_57, ZN => lbl2_sdb_n_123);
  lbl2_sdb_g8632 : AN4D1BWP7T port map(A1 => lbl2_sdb_n_89, A2 => lbl2_sdb_n_78, A3 => lbl2_sdb_n_61, A4 => lbl2_sdb_n_8, Z => lbl2_sdb_n_129);
  lbl2_sdb_g8633 : OAI222D0BWP7T port map(A1 => lbl2_sdb_n_44, A2 => lbl2_sdb_n_76, B1 => lbl2_sdb_n_30, B2 => lbl2_sdb_n_96, C1 => lbl2_sdb_n_60, C2 => lbl2_sdb_n_42, ZN => lbl2_sdb_n_128);
  lbl2_sdb_g8634 : INVD0BWP7T port map(I => lbl2_sdb_n_120, ZN => lbl2_sdb_n_119);
  lbl2_sdb_g8635 : OR2D1BWP7T port map(A1 => lbl2_sdb_n_103, A2 => lbl2_sdb_n_11, Z => lbl2_sdb_n_117);
  lbl2_sdb_g8636 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_97, A2 => lbl2_v_count(4), ZN => lbl2_sdb_n_122);
  lbl2_sdb_g8637 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_98, A2 => lbl2_sdb_n_12, ZN => lbl2_sdb_n_121);
  lbl2_sdb_g8638 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_98, A2 => lbl2_sdb_n_11, ZN => lbl2_sdb_n_120);
  lbl2_sdb_g8639 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_98, A2 => lbl2_v_count(4), ZN => lbl2_sdb_n_118);
  lbl2_sdb_g8640 : INR2XD0BWP7T port map(A1 => lbl2_sdb_n_103, B1 => lbl2_sdb_n_101, ZN => lbl2_sdb_n_116);
  lbl2_sdb_g8641 : OAI211D1BWP7T port map(A1 => lbl2_sdb_n_28, A2 => lbl2_sdb_n_43, B => lbl2_sdb_n_89, C => lbl2_sdb_n_60, ZN => lbl2_sdb_n_115);
  lbl2_sdb_g8642 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_86, A2 => lbl2_sdb_n_54, B => lbl2_sdb_n_28, ZN => lbl2_sdb_n_114);
  lbl2_sdb_g8643 : AOI221D0BWP7T port map(A1 => lbl2_sdb_n_81, A2 => lbl2_sdb_n_2, B1 => lbl2_sdb_n_33, B2 => lbl2_sdb_n_25, C => lbl2_sdb_n_62, ZN => lbl2_sdb_n_113);
  lbl2_sdb_g8644 : OAI21D0BWP7T port map(A1 => lbl2_sdb_n_93, A2 => FE_DBTN18_lbl2_v_count_2, B => lbl2_sdb_n_18, ZN => lbl2_sdb_n_112);
  lbl2_sdb_g8645 : OAI32D1BWP7T port map(A1 => FE_DBTN21_lbl2_h_count_3, A2 => lbl2_v_count(4), A3 => lbl2_sdb_n_78, B1 => lbl2_sdb_n_35, B2 => lbl2_sdb_n_79, ZN => lbl2_sdb_n_111);
  lbl2_sdb_g8646 : NR2D0BWP7T port map(A1 => lbl2_sdb_n_40, A2 => lbl2_sdb_n_93, ZN => lbl2_sdb_n_105);
  lbl2_sdb_g8647 : OAI21D0BWP7T port map(A1 => lbl2_sdb_n_75, A2 => lbl2_sdb_n_50, B => lbl2_sdb_n_93, ZN => lbl2_sdb_n_104);
  lbl2_sdb_g8648 : NR2D0BWP7T port map(A1 => lbl2_sdb_n_93, A2 => lbl2_sdb_n_57, ZN => lbl2_sdb_n_110);
  lbl2_sdb_g8649 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_86, A2 => lbl2_sdb_n_12, ZN => lbl2_sdb_n_109);
  lbl2_sdb_g8650 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_93, A2 => lbl2_sdb_n_27, ZN => lbl2_sdb_n_108);
  lbl2_sdb_g8651 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_87, A2 => lbl2_sdb_n_77, ZN => lbl2_sdb_n_107);
  lbl2_sdb_g8652 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_93, A2 => lbl2_sdb_n_57, ZN => lbl2_sdb_n_106);
  lbl2_sdb_g8653 : INVD0BWP7T port map(I => lbl2_sdb_n_102, ZN => lbl2_sdb_n_101);
  lbl2_sdb_g8654 : INVD0BWP7T port map(I => lbl2_sdb_n_100, ZN => lbl2_sdb_n_99);
  lbl2_sdb_g8655 : CKND1BWP7T port map(I => lbl2_sdb_n_98, ZN => lbl2_sdb_n_97);
  lbl2_sdb_g8656 : AOI22D0BWP7T port map(A1 => lbl2_sdb_n_26, A2 => FE_DBTN21_lbl2_h_count_3, B1 => lbl2_sdb_n_59, B2 => lbl2_h_count(1), ZN => lbl2_sdb_n_96);
  lbl2_sdb_g8657 : ND3D0BWP7T port map(A1 => lbl2_sdb_n_49, A2 => lbl2_sdb_n_22, A3 => lbl2_sdb_n_93, ZN => lbl2_sdb_n_95);
  lbl2_sdb_g8658 : OAI21D0BWP7T port map(A1 => lbl2_sdb_n_79, A2 => lbl2_sdb_n_15, B => lbl2_sdb_n_61, ZN => lbl2_sdb_n_94);
  lbl2_sdb_g8659 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_86, A2 => lbl2_sdb_n_77, ZN => lbl2_sdb_n_103);
  lbl2_sdb_g8660 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_87, A2 => lbl2_sdb_n_93, ZN => lbl2_sdb_n_102);
  lbl2_sdb_g8661 : MOAI22D0BWP7T port map(A1 => lbl2_sdb_n_83, A2 => lbl2_n_150, B1 => lbl2_sdb_n_83, B2 => lbl2_n_150, ZN => lbl2_sdb_n_100);
  lbl2_sdb_g8662 : OAI211D1BWP7T port map(A1 => lbl2_sdb_n_66, A2 => lbl2_sdb_n_9, B => lbl2_sdb_n_83, C => lbl2_sdb_n_20, ZN => lbl2_sdb_n_98);
  lbl2_sdb_g8663 : INVD1BWP7T port map(I => lbl2_sdb_n_77, ZN => lbl2_sdb_n_93);
  lbl2_sdb_g8664 : AO221D0BWP7T port map(A1 => lbl2_sdb_n_53, A2 => lbl2_sdb_n_2, B1 => lbl2_sdb_n_38, B2 => lbl2_sdb_n_12, C => lbl2_sdb_n_56, Z => lbl2_sdb_n_92);
  lbl2_sdb_g8665 : IND3D1BWP7T port map(A1 => lbl2_n_152, B1 => lbl2_sdb_n_71, B2 => lbl2_sdb_n_45, ZN => lbl2_sdb_n_91);
  lbl2_sdb_g8666 : AOI211XD0BWP7T port map(A1 => lbl2_sdb_n_22, A2 => lbl2_sdb_n_12, B => lbl2_sdb_n_64, C => lbl2_sdb_n_52, ZN => lbl2_sdb_n_90);
  lbl2_sdb_g8667 : INVD0BWP7T port map(I => lbl2_sdb_n_89, ZN => lbl2_sdb_n_88);
  lbl2_sdb_g8668 : INVD1BWP7T port map(I => lbl2_sdb_n_87, ZN => lbl2_sdb_n_86);
  lbl2_sdb_g8669 : AOI221D0BWP7T port map(A1 => lbl2_sdb_n_52, A2 => lbl2_v_count(2), B1 => lbl2_sdb_n_55, B2 => lbl2_sdb_n_25, C => lbl2_sdb_n_56, ZN => lbl2_sdb_n_85);
  lbl2_sdb_g8671 : OAI211D1BWP7T port map(A1 => lbl2_sdb_n_58, A2 => lbl2_sdb_n_9, B => lbl2_sdb_n_68, C => lbl2_sdb_n_20, ZN => lbl2_sdb_n_89);
  lbl2_sdb_g8672 : MAOI22D0BWP7T port map(A1 => lbl2_sdb_n_2, A2 => lbl2_sdb_n_66, B1 => lbl2_sdb_n_2, B2 => lbl2_sdb_n_66, ZN => lbl2_sdb_n_87);
  lbl2_sdb_g8673 : IOA21D1BWP7T port map(A1 => lbl2_sdb_n_52, A2 => lbl2_sdb_n_12, B => lbl2_sdb_n_36, ZN => lbl2_sdb_n_82);
  lbl2_sdb_g8674 : IAO21D0BWP7T port map(A1 => lbl2_sdb_n_52, A2 => lbl2_sdb_n_53, B => lbl2_v_count(3), ZN => lbl2_sdb_n_81);
  lbl2_sdb_g8675 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_38, A2 => lbl2_sdb_n_54, B => lbl2_sdb_n_39, ZN => lbl2_sdb_n_80);
  lbl2_sdb_g8676 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_22, A2 => lbl2_sdb_n_66, ZN => lbl2_sdb_n_83);
  lbl2_sdb_g8677 : INVD1BWP7T port map(I => lbl2_sdb_n_79, ZN => lbl2_sdb_n_78);
  lbl2_sdb_g8678 : AOI32D1BWP7T port map(A1 => FE_DBTN21_lbl2_h_count_3, A2 => FE_DBTN20_lbl2_h_count_2, A3 => lbl2_h_count(1), B1 => lbl2_sdb_n_59, B2 => FE_DBTN19_lbl2_h_count_1, ZN => lbl2_sdb_n_76);
  lbl2_sdb_g8679 : MAOI22D0BWP7T port map(A1 => lbl2_sdb_n_51, A2 => lbl2_sdb_n_2, B1 => lbl2_sdb_n_33, B2 => lbl2_sdb_n_2, ZN => lbl2_sdb_n_75);
  lbl2_sdb_g8680 : AOI211XD0BWP7T port map(A1 => lbl2_sdb_n_24, A2 => lbl2_sdb_n_21, B => lbl2_sdb_n_55, C => lbl2_sdb_n_53, ZN => lbl2_sdb_n_74);
  lbl2_sdb_g8681 : OAI22D0BWP7T port map(A1 => lbl2_sdb_n_2, A2 => lbl2_sdb_n_58, B1 => lbl2_n_148, B2 => lbl2_sdb_n_59, ZN => lbl2_sdb_n_79);
  lbl2_sdb_g8682 : MAOI22D0BWP7T port map(A1 => lbl2_sdb_n_26, A2 => lbl2_h_count(3), B1 => lbl2_sdb_n_26, B2 => lbl2_h_count(3), ZN => lbl2_sdb_n_77);
  lbl2_sdb_g8683 : INVD0BWP7T port map(I => lbl2_sdb_n_72, ZN => lbl2_sdb_n_73);
  lbl2_sdb_g8685 : ND4D0BWP7T port map(A1 => lbl2_sdb_n_3, A2 => lbl2_sdb_n_13, A3 => lbl2_v_count(8), A4 => lbl2_v_count(7), ZN => lbl2_sdb_n_67);
  lbl2_sdb_g8686 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_57, A2 => lbl2_v_count(2), ZN => lbl2_sdb_n_72);
  lbl2_sdb_g8687 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_30, A2 => lbl2_sdb_n_60, ZN => lbl2_sdb_n_71);
  lbl2_sdb_g8688 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_57, A2 => lbl2_sdb_n_23, ZN => lbl2_sdb_n_70);
  lbl2_sdb_g8689 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_22, A2 => lbl2_sdb_n_58, ZN => lbl2_sdb_n_68);
  lbl2_sdb_g8690 : OAI32D1BWP7T port map(A1 => FE_DBTN18_lbl2_v_count_2, A2 => lbl2_sdb_n_23, A3 => lbl2_sdb_n_21, B1 => lbl2_n_148, B2 => lbl2_sdb_n_40, ZN => lbl2_sdb_n_65);
  lbl2_sdb_g8691 : OA21D0BWP7T port map(A1 => lbl2_sdb_n_33, A2 => lbl2_sdb_n_19, B => lbl2_sdb_n_49, Z => lbl2_sdb_n_64);
  lbl2_sdb_g8692 : AOI22D0BWP7T port map(A1 => lbl2_sdb_n_0, A2 => lbl2_sdb_n_10, B1 => lbl2_sdb_n_41, B2 => lbl2_h_count(9), ZN => lbl2_sdb_n_63);
  lbl2_sdb_g8693 : MOAI22D0BWP7T port map(A1 => lbl2_sdb_n_36, A2 => lbl2_sdb_n_25, B1 => lbl2_sdb_n_37, B2 => lbl2_n_149, ZN => lbl2_sdb_n_62);
  lbl2_sdb_g8694 : AOI21D0BWP7T port map(A1 => lbl2_h_count(1), A2 => lbl2_h_count(3), B => lbl2_sdb_n_59, ZN => lbl2_sdb_n_66);
  lbl2_sdb_g8695 : INVD1BWP7T port map(I => lbl2_sdb_n_61, ZN => lbl2_sdb_n_60);
  lbl2_sdb_g8696 : INVD1BWP7T port map(I => lbl2_sdb_n_59, ZN => lbl2_sdb_n_58);
  lbl2_sdb_g8697 : INVD1BWP7T port map(I => lbl2_sdb_n_27, ZN => lbl2_sdb_n_57);
  lbl2_sdb_g8698 : HA1D0BWP7T port map(A => lbl2_h_count(3), B => lbl2_h_count(2), CO => lbl2_sdb_n_59, S => lbl2_sdb_n_61);
  lbl2_sdb_g8699 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_37, A2 => FE_DBTN18_lbl2_v_count_2, ZN => lbl2_sdb_n_51);
  lbl2_sdb_g8700 : NR2D0BWP7T port map(A1 => lbl2_sdb_n_29, A2 => lbl2_n_149, ZN => lbl2_sdb_n_50);
  lbl2_sdb_g8701 : AN2D0BWP7T port map(A1 => lbl2_sdb_n_33, A2 => lbl2_n_149, Z => lbl2_sdb_n_56);
  lbl2_sdb_g8702 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_36, A2 => lbl2_v_count(3), ZN => lbl2_sdb_n_55);
  lbl2_sdb_g8703 : ND2D0BWP7T port map(A1 => lbl2_sdb_n_35, A2 => lbl2_sdb_n_23, ZN => lbl2_sdb_n_54);
  lbl2_sdb_g8704 : NR2D1BWP7T port map(A1 => lbl2_n_150, A2 => lbl2_sdb_n_35, ZN => lbl2_sdb_n_53);
  lbl2_sdb_g8705 : AN2D1BWP7T port map(A1 => lbl2_sdb_n_38, A2 => lbl2_sdb_n_8, Z => lbl2_sdb_n_52);
  lbl2_sdb_g8706 : INVD0BWP7T port map(I => lbl2_sdb_n_47, ZN => lbl2_sdb_n_48);
  lbl2_sdb_g8708 : CKMUX2D1BWP7T port map(I0 => lbl2_sdb_n_13, I1 => lbl2_sdb_n_17, S => lbl2_n_153, Z => lbl2_sdb_n_45);
  lbl2_sdb_g8709 : MAOI22D0BWP7T port map(A1 => lbl2_sdb_n_12, A2 => lbl2_v_count(1), B1 => lbl2_sdb_n_15, B2 => lbl2_v_count(1), ZN => lbl2_sdb_n_44);
  lbl2_sdb_g8710 : AOI21D0BWP7T port map(A1 => lbl2_sdb_n_11, A2 => lbl2_v_count(4), B => lbl2_h_count(2), ZN => lbl2_sdb_n_43);
  lbl2_sdb_g8711 : MUX2D1BWP7T port map(I0 => lbl2_sdb_n_11, I1 => lbl2_sdb_n_15, S => lbl2_v_count(1), Z => lbl2_sdb_n_42);
  lbl2_sdb_g8712 : IND2D1BWP7T port map(A1 => lbl2_sdb_n_33, B1 => lbl2_sdb_n_29, ZN => lbl2_sdb_n_49);
  lbl2_sdb_g8713 : IND4D0BWP7T port map(A1 => lbl2_v_count(8), B1 => lbl2_v_count(5), B2 => lbl2_v_count(7), B3 => lbl2_v_count(6), ZN => lbl2_sdb_n_47);
  lbl2_sdb_g8714 : AOI31D0BWP7T port map(A1 => lbl2_v_count(8), A2 => lbl2_v_count(5), A3 => lbl2_v_count(6), B => lbl2_v_count(7), ZN => lbl2_sdb_n_46);
  lbl2_sdb_g8715 : INVD0BWP7T port map(I => lbl2_sdb_n_40, ZN => lbl2_sdb_n_39);
  lbl2_sdb_g8716 : INVD1BWP7T port map(I => lbl2_sdb_n_34, ZN => lbl2_sdb_n_35);
  lbl2_sdb_g8717 : INR2D1BWP7T port map(A1 => game_state(1), B1 => lbl2_sdb_n_16, ZN => lbl2_sdb_n_41);
  lbl2_sdb_g8718 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_24, A2 => lbl2_sdb_n_12, ZN => lbl2_sdb_n_40);
  lbl2_sdb_g8719 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_21, A2 => lbl2_sdb_n_3, ZN => lbl2_sdb_n_38);
  lbl2_sdb_g8720 : NR2D1BWP7T port map(A1 => lbl2_n_150, A2 => lbl2_sdb_n_23, ZN => lbl2_sdb_n_37);
  lbl2_sdb_g8721 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_24, A2 => lbl2_v_count(2), ZN => lbl2_sdb_n_36);
  lbl2_sdb_g8722 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_11, A2 => lbl2_sdb_n_8, ZN => lbl2_sdb_n_34);
  lbl2_sdb_g8723 : NR2D1BWP7T port map(A1 => lbl2_n_150, A2 => lbl2_sdb_n_11, ZN => lbl2_sdb_n_33);
  lbl2_sdb_g8725 : IND3D0BWP7T port map(A1 => game_state(1), B1 => game_state(0), B2 => game_state(2), ZN => lbl2_sdb_n_32);
  lbl2_sdb_g8726 : NR3D0BWP7T port map(A1 => game_state(2), A2 => game_state(0), A3 => game_state(1), ZN => lbl2_sdb_n_31);
  lbl2_sdb_g8727 : AOI21D0BWP7T port map(A1 => FE_DBTN18_lbl2_v_count_2, A2 => lbl2_v_count(3), B => lbl2_sdb_n_14, ZN => lbl2_sdb_n_30);
  lbl2_sdb_g8728 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_24, A2 => FE_DBTN18_lbl2_v_count_2, ZN => lbl2_sdb_n_29);
  lbl2_sdb_g8729 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_23, A2 => lbl2_v_count(2), ZN => lbl2_sdb_n_28);
  lbl2_sdb_g8730 : AOI21D0BWP7T port map(A1 => lbl2_h_count(1), A2 => lbl2_h_count(2), B => lbl2_sdb_n_26, ZN => lbl2_sdb_n_27);
  lbl2_sdb_g8732 : INVD1BWP7T port map(I => lbl2_sdb_n_22, ZN => lbl2_sdb_n_21);
  lbl2_sdb_g8733 : INVD0BWP7T port map(I => lbl2_sdb_n_20, ZN => lbl2_sdb_n_19);
  lbl2_sdb_g8734 : NR2XD0BWP7T port map(A1 => lbl2_h_count(1), A2 => lbl2_h_count(2), ZN => lbl2_sdb_n_26);
  lbl2_sdb_g8735 : NR2D1BWP7T port map(A1 => lbl2_sdb_n_2, A2 => lbl2_n_149, ZN => lbl2_sdb_n_25);
  lbl2_sdb_g8736 : NR2D1BWP7T port map(A1 => lbl2_n_150, A2 => lbl2_v_count(4), ZN => lbl2_sdb_n_24);
  lbl2_sdb_g8737 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_8, A2 => lbl2_v_count(3), ZN => lbl2_sdb_n_23);
  lbl2_sdb_g8738 : NR2D1BWP7T port map(A1 => lbl2_n_149, A2 => lbl2_n_148, ZN => lbl2_sdb_n_22);
  lbl2_sdb_g8739 : ND2D1BWP7T port map(A1 => lbl2_n_149, A2 => lbl2_n_148, ZN => lbl2_sdb_n_20);
  lbl2_sdb_g8740 : INVD1BWP7T port map(I => lbl2_sdb_n_12, ZN => lbl2_sdb_n_11);
  lbl2_sdb_g8741 : ND2D1BWP7T port map(A1 => lbl2_sdb_n_2, A2 => lbl2_n_149, ZN => lbl2_sdb_n_18);
  lbl2_sdb_g8742 : INR2D1BWP7T port map(A1 => lbl2_v_count(6), B1 => lbl2_v_count(5), ZN => lbl2_sdb_n_17);
  lbl2_sdb_g8743 : IND2D1BWP7T port map(A1 => game_state(2), B1 => game_state(0), ZN => lbl2_sdb_n_16);
  lbl2_sdb_g8744 : ND2D1BWP7T port map(A1 => lbl2_v_count(2), A2 => lbl2_v_count(3), ZN => lbl2_sdb_n_15);
  lbl2_sdb_g8745 : NR2D1BWP7T port map(A1 => FE_DBTN18_lbl2_v_count_2, A2 => lbl2_v_count(3), ZN => lbl2_sdb_n_14);
  lbl2_sdb_g8746 : INR2D1BWP7T port map(A1 => lbl2_v_count(5), B1 => lbl2_v_count(6), ZN => lbl2_sdb_n_13);
  lbl2_sdb_g8747 : NR2D1BWP7T port map(A1 => lbl2_v_count(3), A2 => lbl2_v_count(2), ZN => lbl2_sdb_n_12);
  lbl2_sdb_g8748 : INVD0BWP7T port map(I => lbl2_h_count(9), ZN => lbl2_sdb_n_10);
  lbl2_sdb_g8749 : INVD0BWP7T port map(I => lbl2_n_149, ZN => lbl2_sdb_n_9);
  lbl2_sdb_g8750 : INVD1BWP7T port map(I => lbl2_v_count(4), ZN => lbl2_sdb_n_8);
  lbl2_sdb_g8756 : INVD0BWP7T port map(I => lbl2_n_150, ZN => lbl2_sdb_n_3);
  lbl2_sdb_g8757 : INVD1BWP7T port map(I => lbl2_n_148, ZN => lbl2_sdb_n_2);
  lbl2_sdb_g2 : MUX2D0BWP7T port map(I0 => lbl2_sdb_n_25, I1 => lbl2_sdb_n_19, S => lbl2_n_153, Z => lbl2_sdb_n_1);
  lbl2_sdb_g8758 : INR3D0BWP7T port map(A1 => game_state(1), B1 => game_state(2), B2 => game_state(0), ZN => lbl2_sdb_n_0);
  lbl2_sdb_g8759 : XNR2D1BWP7T port map(A1 => lbl2_sdb_n_68, A2 => lbl2_n_150, ZN => lbl2_sdb_n_214);
  lbl0_new_state_reg_0 : LNQD1BWP7T port map(D => lbl0_n_413, EN => lbl0_n_431, Q => lbl0_new_state(0));
  lbl0_new_state_reg_1 : LNQD1BWP7T port map(D => lbl0_n_402, EN => lbl0_n_431, Q => lbl0_new_state(1));
  lbl0_new_state_reg_2 : LNQD1BWP7T port map(D => lbl0_n_377, EN => lbl0_n_431, Q => lbl0_new_state(2));
  lbl0_new_state_reg_3 : LNQD1BWP7T port map(D => lbl0_n_433, EN => lbl0_n_431, Q => lbl0_new_state(3));
  lbl0_new_state_reg_4 : LNQD1BWP7T port map(D => lbl0_n_428, EN => lbl0_n_431, Q => lbl0_new_state(4));
  lbl0_g18423 : OAI211D1BWP7T port map(A1 => lbl0_n_142, A2 => lbl0_n_351, B => lbl0_n_434, C => lbl0_n_224, ZN => lbl0_n_445);
  lbl0_g18424 : OAI211D1BWP7T port map(A1 => lbl0_n_140, A2 => lbl0_n_350, B => lbl0_n_434, C => lbl0_n_222, ZN => lbl0_n_444);
  lbl0_g18425 : AOI211XD0BWP7T port map(A1 => lbl0_n_432, A2 => lbl0_n_138, B => lbl0_n_430, C => lbl0_n_449, ZN => lbl0_n_434);
  lbl0_g18427 : IND4D0BWP7T port map(A1 => lbl0_n_339, B1 => lbl0_n_214, B2 => lbl0_n_216, B3 => lbl0_n_427, ZN => lbl0_n_433);
  lbl0_g18428 : NR4D0BWP7T port map(A1 => lbl0_n_425, A2 => lbl0_n_131, A3 => lbl0_border_0, A4 => lbl0_border_1, ZN => lbl0_n_432);
  lbl0_g18429 : OAI211D1BWP7T port map(A1 => lbl0_n_52, A2 => lbl0_n_191, B => lbl0_n_429, C => lbl0_n_222, ZN => lbl0_n_447);
  lbl0_g18430 : IND3D1BWP7T port map(A1 => lbl0_n_430, B1 => lbl0_n_224, B2 => lbl0_n_240, ZN => lbl0_n_448);
  lbl0_g18432 : INVD0BWP7T port map(I => lbl0_n_430, ZN => lbl0_n_429);
  lbl0_g18433 : AOI211D1BWP7T port map(A1 => lbl0_n_403, A2 => position_0(8), B => lbl0_n_426, C => lbl0_n_412, ZN => lbl0_n_430);
  lbl0_g18434 : IND3D0BWP7T port map(A1 => lbl0_n_243, B1 => lbl0_n_340, B2 => lbl0_n_424, ZN => lbl0_n_428);
  lbl0_g18435 : NR4D0BWP7T port map(A1 => lbl0_n_423, A2 => lbl0_n_249, A3 => lbl0_n_322, A4 => lbl0_n_246, ZN => lbl0_n_427);
  lbl0_g18436 : IND4D0BWP7T port map(A1 => lbl0_n_422, B1 => lbl0_n_138, B2 => lbl0_n_398, B3 => lbl0_n_421, ZN => lbl0_n_426);
  lbl0_g18437 : ND4D0BWP7T port map(A1 => lbl0_n_420, A2 => lbl0_n_414, A3 => lbl0_n_401, A4 => lbl0_n_387, ZN => lbl0_n_425);
  lbl0_g18438 : NR3D0BWP7T port map(A1 => lbl0_n_419, A2 => lbl0_n_325, A3 => lbl0_n_281, ZN => lbl0_n_424);
  lbl0_g18439 : OAI221D0BWP7T port map(A1 => lbl0_n_223, A2 => lbl0_n_285, B1 => lbl0_move_0, B2 => lbl0_n_189, C => lbl0_n_418, ZN => lbl0_n_423);
  lbl0_g18440 : OAI21D0BWP7T port map(A1 => lbl0_n_416, A2 => lbl0_n_208, B => lbl0_n_215, ZN => lbl0_d_position_1(9));
  lbl0_g18441 : OAI211D1BWP7T port map(A1 => position_0(9), A2 => lbl0_n_416, B => lbl0_n_133, C => lbl0_n_132, ZN => lbl0_n_422);
  lbl0_g18442 : AOI211XD0BWP7T port map(A1 => lbl0_n_416, A2 => position_0(9), B => lbl0_n_391, C => lbl0_n_381, ZN => lbl0_n_421);
  lbl0_g18443 : MAOI22D0BWP7T port map(A1 => lbl0_n_417, A2 => lbl0_n_416, B1 => lbl0_n_417, B2 => lbl0_n_416, ZN => lbl0_n_420);
  lbl0_g18444 : AN2D0BWP7T port map(A1 => lbl0_n_417, A2 => lbl0_n_206, Z => lbl0_n_443);
  lbl0_g18445 : OAI31D0BWP7T port map(A1 => lbl0_n_94, A2 => lbl0_n_167, A3 => lbl0_n_406, B => lbl0_n_247, ZN => lbl0_n_419);
  lbl0_g18446 : OAI221D0BWP7T port map(A1 => lbl0_n_405, A2 => lbl0_n_316, B1 => lbl0_n_312, B2 => lbl0_n_404, C => lbl0_n_408, ZN => address(9));
  lbl0_g18447 : AOI21D0BWP7T port map(A1 => lbl0_n_530, A2 => lbl0_n_58, B => lbl0_n_415, ZN => lbl0_n_418);
  lbl0_g18448 : OAI221D0BWP7T port map(A1 => lbl0_n_386, A2 => lbl0_n_316, B1 => lbl0_n_312, B2 => lbl0_n_394, C => lbl0_n_407, ZN => address(8));
  lbl0_g18449 : ND2D1BWP7T port map(A1 => lbl0_n_410, A2 => lbl0_n_349, ZN => address(6));
  lbl0_g18451 : OAI221D0BWP7T port map(A1 => lbl0_n_367, A2 => lbl0_n_316, B1 => lbl0_n_334, B2 => lbl0_n_312, C => lbl0_n_409, ZN => address(7));
  lbl0_g18452 : OAI221D0BWP7T port map(A1 => lbl0_n_316, A2 => position_0(5), B1 => position_1(5), B2 => lbl0_n_312, C => lbl0_n_411, ZN => address(5));
  lbl0_g18453 : OAI21D0BWP7T port map(A1 => lbl0_n_403, A2 => lbl0_n_208, B => lbl0_n_158, ZN => lbl0_d_position_1(8));
  lbl0_g18454 : INR3D0BWP7T port map(A1 => lbl0_n_406, B1 => lbl0_n_94, B2 => lbl0_n_167, ZN => lbl0_n_415);
  lbl0_g18455 : MAOI22D0BWP7T port map(A1 => lbl0_n_403, A2 => lbl0_n_397, B1 => lbl0_n_403, B2 => lbl0_n_397, ZN => lbl0_n_414);
  lbl0_g18456 : MOAI22D0BWP7T port map(A1 => lbl0_n_405, A2 => lbl0_next_direction_0(0), B1 => lbl0_next_direction_0(0), B2 => position_0(9), ZN => lbl0_n_417);
  lbl0_g18457 : MAOI22D0BWP7T port map(A1 => lbl0_next_direction_1(0), A2 => position_1(9), B1 => lbl0_n_404, B2 => lbl0_next_direction_1(0), ZN => lbl0_n_416);
  lbl0_g18458 : OR3D0BWP7T port map(A1 => lbl0_n_323, A2 => lbl0_n_281, A3 => lbl0_n_395, Z => lbl0_n_413);
  lbl0_g18459 : NR2XD0BWP7T port map(A1 => lbl0_n_403, A2 => position_0(8), ZN => lbl0_n_412);
  lbl0_g18461 : AO21D0BWP7T port map(A1 => lbl0_n_397, A2 => lbl0_n_206, B => lbl0_n_211, Z => lbl0_d_position_0(8));
  lbl0_g18462 : AOI22D0BWP7T port map(A1 => lbl0_n_400, A2 => position_1(5), B1 => lbl0_n_338, B2 => position_0(5), ZN => lbl0_n_411);
  lbl0_g18463 : AOI22D0BWP7T port map(A1 => lbl0_n_400, A2 => position_1(6), B1 => lbl0_n_338, B2 => position_0(6), ZN => lbl0_n_410);
  lbl0_g18464 : AOI22D0BWP7T port map(A1 => lbl0_n_400, A2 => position_1(7), B1 => lbl0_n_338, B2 => position_0(7), ZN => lbl0_n_409);
  lbl0_g18465 : AOI22D0BWP7T port map(A1 => lbl0_n_400, A2 => position_1(9), B1 => lbl0_n_338, B2 => position_0(9), ZN => lbl0_n_408);
  lbl0_g18466 : AOI22D0BWP7T port map(A1 => lbl0_n_400, A2 => position_1(8), B1 => lbl0_n_338, B2 => position_0(8), ZN => lbl0_n_407);
  lbl0_g18467 : CKAN2D1BWP7T port map(A1 => lbl0_n_399, A2 => read_memory_in(0), Z => lbl0_d_read_data_reg(0));
  lbl0_g18468 : CKAN2D1BWP7T port map(A1 => lbl0_n_399, A2 => read_memory_in(5), Z => lbl0_d_read_data_reg(5));
  lbl0_g18469 : CKAN2D1BWP7T port map(A1 => lbl0_n_399, A2 => read_memory_in(3), Z => lbl0_d_read_data_reg(3));
  lbl0_g18470 : CKAN2D1BWP7T port map(A1 => lbl0_n_399, A2 => read_memory_in(2), Z => lbl0_d_read_data_reg(2));
  lbl0_g18471 : CKAN2D1BWP7T port map(A1 => lbl0_n_399, A2 => read_memory_in(1), Z => lbl0_d_read_data_reg(1));
  lbl0_g18472 : CKAN2D1BWP7T port map(A1 => lbl0_n_399, A2 => read_memory_in(4), Z => lbl0_d_read_data_reg(4));
  lbl0_g18473 : CKAN2D1BWP7T port map(A1 => lbl0_n_399, A2 => read_memory_in(6), Z => lbl0_d_read_data_reg(6));
  lbl0_g18474 : IND4D0BWP7T port map(A1 => lbl0_n_382, B1 => lbl0_n_209, B2 => lbl0_n_340, B3 => lbl0_n_356, ZN => lbl0_n_402);
  lbl0_g18475 : NR4D0BWP7T port map(A1 => lbl0_n_396, A2 => lbl0_n_359, A3 => lbl0_n_363, A4 => lbl0_n_362, ZN => lbl0_n_401);
  lbl0_g18476 : CKAN2D1BWP7T port map(A1 => lbl0_n_399, A2 => read_memory_in(7), Z => lbl0_d_read_data_reg(7));
  lbl0_g18477 : NR4D0BWP7T port map(A1 => lbl0_n_390, A2 => lbl0_n_353, A3 => lbl0_busy_count(6), A4 => lbl0_busy_count(5), ZN => lbl0_n_406);
  lbl0_g18478 : MAOI22D0BWP7T port map(A1 => lbl0_n_393, A2 => position_0(9), B1 => lbl0_n_393, B2 => position_0(9), ZN => lbl0_n_405);
  lbl0_g18479 : MAOI22D0BWP7T port map(A1 => lbl0_n_392, A2 => lbl0_n_204, B1 => lbl0_n_392, B2 => lbl0_n_204, ZN => lbl0_n_404);
  lbl0_g18480 : MAOI22D0BWP7T port map(A1 => lbl0_next_direction_1(0), A2 => position_1(8), B1 => lbl0_n_394, B2 => lbl0_next_direction_1(0), ZN => lbl0_n_403);
  lbl0_g18481 : NR4D0BWP7T port map(A1 => lbl0_n_380, A2 => lbl0_n_388, A3 => lbl0_n_298, A4 => lbl0_n_233, ZN => lbl0_n_398);
  lbl0_g18483 : NR4D0BWP7T port map(A1 => lbl0_n_374, A2 => lbl0_n_338, A3 => lbl0_n_311, A4 => lbl0_n_267, ZN => lbl0_n_400);
  lbl0_g18484 : AN4D1BWP7T port map(A1 => lbl0_n_375, A2 => lbl0_n_268, A3 => lbl0_n_141, A4 => lbl0_n_140, Z => lbl0_n_399);
  lbl0_g18485 : MOAI22D0BWP7T port map(A1 => lbl0_n_384, A2 => lbl0_n_366, B1 => lbl0_n_384, B2 => lbl0_n_366, ZN => lbl0_n_396);
  lbl0_g18486 : AO21D0BWP7T port map(A1 => lbl0_n_385, A2 => lbl0_n_206, B => lbl0_n_211, Z => lbl0_d_position_0(7));
  lbl0_g18487 : OAI211D0BWP7T port map(A1 => lbl0_move_1, A2 => lbl0_n_216, B => lbl0_n_389, C => lbl0_n_299, ZN => lbl0_n_395);
  lbl0_g18488 : MOAI22D0BWP7T port map(A1 => lbl0_n_386, A2 => lbl0_next_direction_0(0), B1 => lbl0_next_direction_0(0), B2 => position_0(8), ZN => lbl0_n_397);
  lbl0_g18489 : MAOI22D0BWP7T port map(A1 => lbl0_n_348, A2 => lbl0_n_90, B1 => lbl0_n_369, B2 => lbl0_n_90, ZN => lbl0_n_394);
  lbl0_g18490 : NR2D0BWP7T port map(A1 => lbl0_n_383, A2 => lbl0_state(1), ZN => lbl0_n_431);
  lbl0_g18491 : MAOI22D0BWP7T port map(A1 => lbl0_n_376, A2 => lbl0_n_114, B1 => lbl0_n_376, B2 => lbl0_n_114, ZN => lbl0_n_393);
  lbl0_g18492 : AOI22D0BWP7T port map(A1 => lbl0_n_357, A2 => lbl0_n_91, B1 => lbl0_n_306, B2 => position_1(8), ZN => lbl0_n_392);
  lbl0_g18493 : OAI221D0BWP7T port map(A1 => lbl0_n_331, A2 => position_0(6), B1 => position_0(5), B2 => lbl0_n_137, C => lbl0_n_378, ZN => lbl0_n_391);
  lbl0_g18494 : AOI21D0BWP7T port map(A1 => lbl0_n_370, A2 => lbl0_n_2, B => test_button, ZN => lbl0_n_390);
  lbl0_g18495 : NR2D0BWP7T port map(A1 => lbl0_n_373, A2 => lbl0_n_339, ZN => lbl0_n_389);
  lbl0_g18496 : OAI221D0BWP7T port map(A1 => lbl0_n_257, A2 => position_1(1), B1 => position_1(0), B2 => lbl0_n_135, C => lbl0_n_379, ZN => lbl0_n_388);
  lbl0_g18497 : NR4D0BWP7T port map(A1 => lbl0_n_345, A2 => lbl0_n_352, A3 => lbl0_n_302, A4 => lbl0_n_301, ZN => lbl0_n_387);
  lbl0_g18498 : INVD0BWP7T port map(I => lbl0_n_384, ZN => lbl0_n_385);
  lbl0_g18499 : IIND4D0BWP7T port map(A1 => lbl0_n_295, A2 => lbl0_n_455, B1 => lbl0_n_358, B2 => lbl0_n_279, ZN => lbl0_n_383);
  lbl0_g18500 : IND4D0BWP7T port map(A1 => lbl0_n_322, B1 => lbl0_n_261, B2 => lbl0_n_276, B3 => lbl0_n_354, ZN => lbl0_n_382);
  lbl0_g18501 : OAI21D0BWP7T port map(A1 => lbl0_n_365, A2 => lbl0_n_208, B => lbl0_n_158, ZN => lbl0_d_position_1(7));
  lbl0_g18502 : MOAI22D0BWP7T port map(A1 => lbl0_n_366, A2 => lbl0_n_61, B1 => lbl0_n_366, B2 => lbl0_n_61, ZN => lbl0_n_381);
  lbl0_g18503 : MAOI22D0BWP7T port map(A1 => lbl0_n_368, A2 => position_0(8), B1 => lbl0_n_368, B2 => position_0(8), ZN => lbl0_n_386);
  lbl0_g18504 : MAOI22D0BWP7T port map(A1 => lbl0_next_direction_0(0), A2 => position_0(7), B1 => lbl0_n_367, B2 => lbl0_next_direction_0(0), ZN => lbl0_n_384);
  lbl0_g18505 : OAI221D0BWP7T port map(A1 => lbl0_n_314, A2 => position_0(2), B1 => position_0(0), B2 => lbl0_n_237, C => lbl0_n_371, ZN => lbl0_n_380);
  lbl0_g18506 : AOI221D0BWP7T port map(A1 => lbl0_n_257, A2 => position_1(1), B1 => lbl0_n_135, B2 => position_1(0), C => lbl0_n_360, ZN => lbl0_n_379);
  lbl0_g18507 : AOI221D0BWP7T port map(A1 => lbl0_n_331, A2 => position_0(6), B1 => lbl0_n_137, B2 => position_0(5), C => lbl0_n_364, ZN => lbl0_n_378);
  lbl0_g18508 : ND2D0BWP7T port map(A1 => lbl0_n_372, A2 => lbl0_n_356, ZN => lbl0_n_377);
  lbl0_g18509 : INVD0BWP7T port map(I => lbl0_n_374, ZN => lbl0_n_375);
  lbl0_g18510 : ND4D0BWP7T port map(A1 => lbl0_n_327, A2 => lbl0_n_297, A3 => lbl0_n_274, A4 => lbl0_n_245, ZN => lbl0_n_373);
  lbl0_g18511 : OAI221D0BWP7T port map(A1 => lbl0_n_305, A2 => lbl0_n_286, B1 => lbl0_n_68, B2 => lbl0_n_277, C => lbl0_n_361, ZN => address(4));
  lbl0_g18512 : AOI22D0BWP7T port map(A1 => lbl0_n_355, A2 => lbl0_n_114, B1 => lbl0_n_309, B2 => position_0(8), ZN => lbl0_n_376);
  lbl0_g18513 : ND3D0BWP7T port map(A1 => lbl0_n_358, A2 => lbl0_n_213, A3 => lbl0_n_101, ZN => lbl0_n_374);
  lbl0_g18514 : NR3D0BWP7T port map(A1 => lbl0_n_336, A2 => lbl0_n_323, A3 => lbl0_n_246, ZN => lbl0_n_372);
  lbl0_g18515 : AOI221D0BWP7T port map(A1 => lbl0_n_314, A2 => position_0(2), B1 => lbl0_n_237, B2 => position_0(0), C => lbl0_n_347, ZN => lbl0_n_371);
  lbl0_g18516 : OAI221D0BWP7T port map(A1 => lbl0_n_307, A2 => lbl0_n_286, B1 => lbl0_n_83, B2 => lbl0_n_277, C => lbl0_n_346, ZN => address(3));
  lbl0_g18517 : OAI221D0BWP7T port map(A1 => lbl0_n_319, A2 => lbl0_n_286, B1 => lbl0_n_80, B2 => lbl0_n_277, C => lbl0_n_343, ZN => address(2));
  lbl0_g18518 : MAOI222D0BWP7T port map(A => lbl0_busy_count(3), B => lbl0_n_502, C => lbl0_n_308, ZN => lbl0_n_370);
  lbl0_g18519 : OAI222D0BWP7T port map(A1 => lbl0_n_318, A2 => lbl0_n_73, B1 => lbl0_n_241, B2 => lbl0_n_289, C1 => lbl0_n_239, C2 => lbl0_n_54, ZN => write_memory(4));
  lbl0_g18520 : OA21D0BWP7T port map(A1 => lbl0_n_341, A2 => lbl0_n_64, B => lbl0_n_357, Z => lbl0_n_369);
  lbl0_g18521 : AO21D0BWP7T port map(A1 => lbl0_n_332, A2 => lbl0_n_206, B => lbl0_n_211, Z => lbl0_d_position_0(6));
  lbl0_g18522 : OAI21D0BWP7T port map(A1 => lbl0_n_331, A2 => lbl0_n_208, B => lbl0_n_210, ZN => lbl0_d_position_1(6));
  lbl0_g18523 : AO222D0BWP7T port map(A1 => lbl0_n_320, A2 => lbl0_read_data_reg(2), B1 => lbl0_n_293, B2 => lbl0_n_147, C1 => lbl0_n_291, C2 => lbl0_n_150, Z => write_memory(2));
  lbl0_g18524 : INVD0BWP7T port map(I => lbl0_n_366, ZN => lbl0_n_365);
  lbl0_g18525 : MOAI22D0BWP7T port map(A1 => lbl0_n_330, A2 => lbl0_n_68, B1 => lbl0_n_330, B2 => lbl0_n_68, ZN => lbl0_n_364);
  lbl0_g18526 : MOAI22D0BWP7T port map(A1 => lbl0_n_331, A2 => lbl0_n_332, B1 => lbl0_n_137, B2 => lbl0_n_136, ZN => lbl0_n_363);
  lbl0_g18527 : MOAI22D0BWP7T port map(A1 => lbl0_n_137, A2 => lbl0_n_136, B1 => lbl0_n_331, B2 => lbl0_n_332, ZN => lbl0_n_362);
  lbl0_g18528 : OAI22D0BWP7T port map(A1 => lbl0_n_329, A2 => lbl0_n_208, B1 => lbl0_n_158, B2 => start_position_0(3), ZN => lbl0_d_position_1(4));
  lbl0_g18529 : AOI22D0BWP7T port map(A1 => lbl0_n_330, A2 => lbl0_n_287, B1 => lbl0_n_278, B2 => position_1(4), ZN => lbl0_n_361);
  lbl0_g18531 : MOAI22D0BWP7T port map(A1 => lbl0_n_333, A2 => position_1(6), B1 => lbl0_n_333, B2 => position_1(6), ZN => lbl0_n_360);
  lbl0_g18532 : MOAI22D0BWP7T port map(A1 => lbl0_n_330, A2 => lbl0_n_305, B1 => lbl0_n_330, B2 => lbl0_n_305, ZN => lbl0_n_359);
  lbl0_g18533 : AOI22D0BWP7T port map(A1 => lbl0_n_342, A2 => lbl0_n_114, B1 => lbl0_n_309, B2 => lbl0_n_113, ZN => lbl0_n_368);
  lbl0_g18534 : MAOI22D0BWP7T port map(A1 => lbl0_n_335, A2 => lbl0_n_114, B1 => lbl0_n_335, B2 => lbl0_n_114, ZN => lbl0_n_367);
  lbl0_g18535 : MOAI22D0BWP7T port map(A1 => lbl0_n_334, A2 => lbl0_next_direction_1(0), B1 => lbl0_next_direction_1(0), B2 => position_1(7), ZN => lbl0_n_366);
  lbl0_g18536 : IND2D0BWP7T port map(A1 => position_0(8), B1 => lbl0_n_342, ZN => lbl0_n_355);
  lbl0_g18537 : OAI221D0BWP7T port map(A1 => lbl0_n_277, A2 => lbl0_n_82, B1 => lbl0_n_135, B2 => lbl0_n_286, C => lbl0_n_324, ZN => address(0));
  lbl0_g18538 : OAI221D0BWP7T port map(A1 => lbl0_n_257, A2 => lbl0_n_286, B1 => lbl0_n_84, B2 => lbl0_n_277, C => lbl0_n_328, ZN => address(1));
  lbl0_g18539 : AO21D0BWP7T port map(A1 => lbl0_n_320, A2 => lbl0_read_data_reg(0), B => lbl0_n_326, Z => write_memory(0));
  lbl0_g18540 : OAI21D0BWP7T port map(A1 => lbl0_n_318, A2 => lbl0_n_75, B => lbl0_n_289, ZN => write_memory(7));
  lbl0_g18541 : AO21D0BWP7T port map(A1 => lbl0_n_320, A2 => lbl0_read_data_reg(3), B => lbl0_n_291, Z => write_memory(3));
  lbl0_g18542 : OAI21D0BWP7T port map(A1 => lbl0_n_319, A2 => lbl0_n_207, B => lbl0_n_215, ZN => lbl0_d_position_0(2));
  lbl0_g18543 : AOI211D0BWP7T port map(A1 => lbl0_n_284, A2 => lbl0_n_532, B => lbl0_n_300, C => lbl0_n_231, ZN => lbl0_n_354);
  lbl0_g18544 : AN3D0BWP7T port map(A1 => lbl0_n_308, A2 => lbl0_busy_count(3), A3 => lbl0_busy_count(4), Z => lbl0_n_353);
  lbl0_g18545 : OAI21D0BWP7T port map(A1 => lbl0_n_314, A2 => lbl0_n_208, B => lbl0_n_158, ZN => lbl0_d_position_1(2));
  lbl0_g18546 : NR4D0BWP7T port map(A1 => lbl0_n_272, A2 => lbl0_n_535, A3 => lbl0_n_121, A4 => lbl0_n_100, ZN => lbl0_n_358);
  lbl0_g18547 : ND2D1BWP7T port map(A1 => lbl0_n_341, A2 => lbl0_n_64, ZN => lbl0_n_357);
  lbl0_g18548 : AN3D0BWP7T port map(A1 => lbl0_n_337, A2 => lbl0_n_245, A3 => lbl0_n_179, Z => lbl0_n_356);
  lbl0_g18549 : CKXOR2D0BWP7T port map(A1 => lbl0_n_319, A2 => lbl0_n_314, Z => lbl0_n_352);
  lbl0_g18550 : OAI222D0BWP7T port map(A1 => lbl0_n_318, A2 => lbl0_n_74, B1 => lbl0_n_199, B2 => lbl0_n_54, C1 => lbl0_n_197, C2 => lbl0_n_289, ZN => write_memory(5));
  lbl0_g18551 : AOI32D1BWP7T port map(A1 => lbl0_n_296, A2 => lbl0_n_285, A3 => lbl0_n_65, B1 => lbl0_n_310, B2 => lbl0_next_layer_0, ZN => lbl0_n_351);
  lbl0_g18552 : AOI32D1BWP7T port map(A1 => lbl0_n_296, A2 => lbl0_n_285, A3 => lbl0_n_81, B1 => lbl0_n_310, B2 => lbl0_next_layer_1, ZN => lbl0_n_350);
  lbl0_g18553 : AOI22D0BWP7T port map(A1 => lbl0_n_311, A2 => lbl0_n_259, B1 => lbl0_n_315, B2 => lbl0_n_260, ZN => lbl0_n_349);
  lbl0_g18554 : MOAI22D0BWP7T port map(A1 => lbl0_n_303, A2 => lbl0_n_208, B1 => lbl0_n_157, B2 => start_position_1(3), ZN => lbl0_d_position_1(3));
  lbl0_g18555 : MOAI22D0BWP7T port map(A1 => lbl0_n_307, A2 => lbl0_n_207, B1 => lbl0_n_157, B2 => start_position_0(3), ZN => lbl0_d_position_0(3));
  lbl0_g18556 : MOAI22D0BWP7T port map(A1 => lbl0_n_306, A2 => lbl0_n_64, B1 => lbl0_n_306, B2 => lbl0_n_64, ZN => lbl0_n_348);
  lbl0_g18557 : MOAI22D0BWP7T port map(A1 => lbl0_n_304, A2 => lbl0_n_83, B1 => lbl0_n_304, B2 => lbl0_n_83, ZN => lbl0_n_347);
  lbl0_g18558 : AOI22D0BWP7T port map(A1 => lbl0_n_304, A2 => lbl0_n_287, B1 => lbl0_n_278, B2 => position_1(3), ZN => lbl0_n_346);
  lbl0_g18559 : MOAI22D0BWP7T port map(A1 => lbl0_n_304, A2 => lbl0_n_307, B1 => lbl0_n_304, B2 => lbl0_n_307, ZN => lbl0_n_345);
  lbl0_g18561 : AOI22D0BWP7T port map(A1 => lbl0_n_313, A2 => lbl0_n_287, B1 => lbl0_n_278, B2 => position_1(2), ZN => lbl0_n_343);
  lbl0_g18562 : AO222D0BWP7T port map(A1 => lbl0_n_320, A2 => lbl0_read_data_reg(1), B1 => lbl0_n_293, B2 => lbl0_n_198, C1 => lbl0_n_291, C2 => lbl0_n_196, Z => write_memory(1));
  lbl0_g18563 : NR3D0BWP7T port map(A1 => lbl0_n_295, A2 => lbl0_n_213, A3 => lbl0_busy_count(4), ZN => pulse_audio);
  lbl0_g18564 : MOAI22D0BWP7T port map(A1 => lbl0_n_263, A2 => position_1(10), B1 => lbl0_n_283, B2 => position_1(10), ZN => lbl0_n_499);
  lbl0_g18565 : NR2D1BWP7T port map(A1 => lbl0_n_305, A2 => lbl0_n_207, ZN => lbl0_n_441);
  lbl0_g18566 : IND3D0BWP7T port map(A1 => lbl0_n_214, B1 => lbl0_n_56, B2 => lbl0_n_284, ZN => lbl0_n_337);
  lbl0_g18567 : ND3D0BWP7T port map(A1 => lbl0_n_275, A2 => lbl0_n_321, A3 => lbl0_n_247, ZN => lbl0_n_336);
  lbl0_g18568 : NR2XD0BWP7T port map(A1 => lbl0_n_309, A2 => position_0(7), ZN => lbl0_n_342);
  lbl0_g18569 : NR2XD0BWP7T port map(A1 => lbl0_n_306, A2 => position_1(7), ZN => lbl0_n_341);
  lbl0_g18570 : INR2D0BWP7T port map(A1 => lbl0_n_321, B1 => lbl0_n_242, ZN => lbl0_n_340);
  lbl0_g18571 : OAI222D0BWP7T port map(A1 => lbl0_n_179, A2 => lbl0_state(2), B1 => lbl0_n_285, B2 => lbl0_n_218, C1 => lbl0_n_106, C2 => lbl0_n_164, ZN => lbl0_n_339);
  lbl0_g18572 : OAI21D0BWP7T port map(A1 => lbl0_n_286, A2 => lbl0_n_76, B => lbl0_n_277, ZN => lbl0_n_338);
  lbl0_g18573 : INVD0BWP7T port map(I => lbl0_n_333, ZN => lbl0_n_332);
  lbl0_g18574 : INVD0BWP7T port map(I => lbl0_n_330, ZN => lbl0_n_329);
  lbl0_g18575 : AOI22D0BWP7T port map(A1 => lbl0_n_256, A2 => lbl0_n_287, B1 => lbl0_n_278, B2 => position_1(1), ZN => lbl0_n_328);
  lbl0_g18576 : AOI22D0BWP7T port map(A1 => lbl0_n_279, A2 => lbl0_n_212, B1 => lbl0_n_166, B2 => lbl0_state(0), ZN => lbl0_n_327);
  lbl0_g18577 : OAI22D0BWP7T port map(A1 => lbl0_n_294, A2 => lbl0_n_239, B1 => lbl0_n_290, B2 => lbl0_n_241, ZN => lbl0_n_326);
  lbl0_g18578 : OAI22D0BWP7T port map(A1 => lbl0_n_273, A2 => lbl0_n_284, B1 => lbl0_n_279, B2 => lbl0_n_213, ZN => lbl0_n_325);
  lbl0_g18579 : AOI22D0BWP7T port map(A1 => lbl0_n_287, A2 => lbl0_n_236, B1 => lbl0_n_278, B2 => position_1(0), ZN => lbl0_n_324);
  lbl0_g18580 : MOAI22D0BWP7T port map(A1 => lbl0_n_194, A2 => lbl0_n_61, B1 => lbl0_n_194, B2 => lbl0_n_61, ZN => lbl0_n_335);
  lbl0_g18581 : MAOI22D0BWP7T port map(A1 => lbl0_n_203, A2 => lbl0_n_193, B1 => lbl0_n_203, B2 => lbl0_n_193, ZN => lbl0_n_334);
  lbl0_g18582 : AOI22D0BWP7T port map(A1 => lbl0_n_260, A2 => lbl0_n_76, B1 => lbl0_next_direction_0(0), B2 => position_0(6), ZN => lbl0_n_333);
  lbl0_g18583 : AOI22D0BWP7T port map(A1 => lbl0_n_259, A2 => lbl0_n_55, B1 => lbl0_next_direction_1(0), B2 => position_1(6), ZN => lbl0_n_331);
  lbl0_g18584 : MOAI22D0BWP7T port map(A1 => lbl0_n_280, A2 => position_1(4), B1 => lbl0_n_280, B2 => position_1(4), ZN => lbl0_n_330);
  lbl0_g18585 : INVD0BWP7T port map(I => lbl0_n_317, ZN => lbl0_n_318);
  lbl0_g18586 : INVD1BWP7T port map(I => lbl0_n_315, ZN => lbl0_n_316);
  lbl0_g18587 : INVD0BWP7T port map(I => lbl0_n_314, ZN => lbl0_n_313);
  lbl0_g18588 : INVD0BWP7T port map(I => lbl0_n_312, ZN => lbl0_n_311);
  lbl0_g18589 : MOAI22D0BWP7T port map(A1 => lbl0_n_265, A2 => position_0(10), B1 => lbl0_n_264, B2 => position_0(10), ZN => lbl0_n_498);
  lbl0_g18590 : OAI222D0BWP7T port map(A1 => lbl0_n_228, A2 => position_1(10), B1 => FE_DBTN22_position_1_10, B2 => lbl0_n_229, C1 => lbl0_next_direction_1(0), C2 => lbl0_n_205, ZN => lbl0_n_497);
  lbl0_g18591 : OAI21D0BWP7T port map(A1 => lbl0_n_255, A2 => lbl0_n_208, B => lbl0_n_215, ZN => lbl0_d_position_1(1));
  lbl0_g18592 : OAI21D0BWP7T port map(A1 => lbl0_n_251, A2 => position_0(10), B => lbl0_n_282, ZN => lbl0_n_500);
  lbl0_g18593 : NR3D0BWP7T port map(A1 => lbl0_n_216, A2 => lbl0_n_285, A3 => lbl0_state(1), ZN => lbl0_n_323);
  lbl0_g18594 : INR2D0BWP7T port map(A1 => lbl0_n_221, B1 => lbl0_n_285, ZN => lbl0_n_322);
  lbl0_g18595 : IND2D0BWP7T port map(A1 => lbl0_n_223, B1 => lbl0_n_285, ZN => lbl0_n_321);
  lbl0_g18596 : ND2D1BWP7T port map(A1 => lbl0_n_54, A2 => lbl0_n_289, ZN => lbl0_n_320);
  lbl0_g18597 : AOI211XD0BWP7T port map(A1 => lbl0_n_235, A2 => position_0(2), B => lbl0_n_190, C => lbl0_n_186, ZN => lbl0_n_319);
  lbl0_g18598 : ND2D1BWP7T port map(A1 => lbl0_n_290, A2 => lbl0_n_294, ZN => lbl0_n_317);
  lbl0_g18599 : NR2XD0BWP7T port map(A1 => lbl0_n_286, A2 => lbl0_next_direction_0(0), ZN => lbl0_n_315);
  lbl0_g18600 : AOI211XD0BWP7T port map(A1 => lbl0_n_234, A2 => position_1(2), B => lbl0_n_53, C => lbl0_n_51, ZN => lbl0_n_314);
  lbl0_g18601 : ND2D1BWP7T port map(A1 => lbl0_n_287, A2 => lbl0_n_55, ZN => lbl0_n_312);
  lbl0_g18602 : INVD0BWP7T port map(I => lbl0_n_304, ZN => lbl0_n_303);
  lbl0_g18603 : MOAI22D0BWP7T port map(A1 => lbl0_n_256, A2 => lbl0_n_257, B1 => lbl0_n_236, B2 => lbl0_n_135, ZN => lbl0_n_302);
  lbl0_g18604 : MOAI22D0BWP7T port map(A1 => lbl0_n_236, A2 => lbl0_n_135, B1 => lbl0_n_256, B2 => lbl0_n_257, ZN => lbl0_n_301);
  lbl0_g18605 : OAI21D0BWP7T port map(A1 => lbl0_n_257, A2 => lbl0_n_207, B => lbl0_n_215, ZN => lbl0_d_position_0(1));
  lbl0_g18606 : IAO21D0BWP7T port map(A1 => lbl0_n_249, A2 => lbl0_n_536, B => lbl0_n_284, ZN => lbl0_n_300);
  lbl0_g18607 : IND3D0BWP7T port map(A1 => lbl0_n_214, B1 => lbl0_move_0, B2 => lbl0_n_285, ZN => lbl0_n_299);
  lbl0_g18608 : OAI22D0BWP7T port map(A1 => lbl0_n_256, A2 => lbl0_n_84, B1 => lbl0_n_255, B2 => position_0(1), ZN => lbl0_n_298);
  lbl0_g18609 : AOI22D0BWP7T port map(A1 => lbl0_n_262, A2 => start_between, B1 => lbl0_n_161, B2 => lbl0_n_5, ZN => lbl0_n_297);
  lbl0_g18610 : INR3D0BWP7T port map(A1 => lbl0_n_268, B1 => lbl0_n_180, B2 => lbl0_n_284, ZN => lbl0_n_310);
  lbl0_g18611 : AOI21D0BWP7T port map(A1 => lbl0_n_113, A2 => lbl0_n_61, B => lbl0_n_194, ZN => lbl0_n_309);
  lbl0_g18612 : OAI22D0BWP7T port map(A1 => lbl0_n_250, A2 => test_button, B1 => lbl0_n_437, B2 => lbl0_n_4, ZN => lbl0_n_308);
  lbl0_g18613 : AOI22D0BWP7T port map(A1 => lbl0_n_253, A2 => position_0(3), B1 => lbl0_n_230, B2 => lbl0_n_83, ZN => lbl0_n_307);
  lbl0_g18614 : IAO21D0BWP7T port map(A1 => lbl0_n_91, A2 => position_1(7), B => lbl0_n_193, ZN => lbl0_n_306);
  lbl0_g18615 : MAOI22D0BWP7T port map(A1 => lbl0_n_258, A2 => lbl0_n_68, B1 => lbl0_n_258, B2 => lbl0_n_68, ZN => lbl0_n_305);
  lbl0_g18616 : MOAI22D0BWP7T port map(A1 => lbl0_n_269, A2 => position_1(3), B1 => lbl0_n_269, B2 => position_1(3), ZN => lbl0_n_304);
  lbl0_g18617 : INVD0BWP7T port map(I => lbl0_n_293, ZN => lbl0_n_294);
  lbl0_g18618 : INVD0BWP7T port map(I => lbl0_n_54, ZN => lbl0_n_292);
  lbl0_g18619 : INVD0BWP7T port map(I => lbl0_n_291, ZN => lbl0_n_290);
  lbl0_g18620 : INVD1BWP7T port map(I => lbl0_n_288, ZN => lbl0_n_289);
  lbl0_g18621 : INVD1BWP7T port map(I => lbl0_n_285, ZN => lbl0_n_284);
  lbl0_g18622 : OAI221D0BWP7T port map(A1 => ramps(5), A2 => lbl0_n_99, B1 => lbl0_n_95, B2 => ramps(7), C => lbl0_n_252, ZN => lbl0_n_283);
  lbl0_g18623 : OAI21D0BWP7T port map(A1 => lbl0_n_183, A2 => lbl0_n_232, B => position_0(10), ZN => lbl0_n_282);
  lbl0_g18624 : INR2D1BWP7T port map(A1 => lbl0_n_268, B1 => lbl0_n_187, ZN => lbl0_n_296);
  lbl0_g18625 : INR3D0BWP7T port map(A1 => lbl0_n_439, B1 => lbl0_busy_count(5), B2 => lbl0_busy_count(6), ZN => lbl0_n_295);
  lbl0_g18626 : NR2D1BWP7T port map(A1 => lbl0_n_270, A2 => position_0(10), ZN => lbl0_n_293);
  lbl0_g18628 : NR2D1BWP7T port map(A1 => lbl0_n_271, A2 => position_1(10), ZN => lbl0_n_291);
  lbl0_g18629 : NR2D1BWP7T port map(A1 => lbl0_n_271, A2 => FE_DBTN22_position_1_10, ZN => lbl0_n_288);
  lbl0_g18630 : NR2D1BWP7T port map(A1 => lbl0_n_267, A2 => lbl0_n_140, ZN => lbl0_n_287);
  lbl0_g18631 : OR2D1BWP7T port map(A1 => lbl0_n_267, A2 => lbl0_n_142, Z => lbl0_n_286);
  lbl0_g18632 : OAI221D1BWP7T port map(A1 => lbl0_n_126, A2 => lbl0_n_79, B1 => lbl0_mem_com_state(2), B2 => lbl0_n_123, C => lbl0_n_128, ZN => lbl0_n_285);
  lbl0_g18633 : OAI21D0BWP7T port map(A1 => lbl0_n_208, A2 => lbl0_n_237, B => lbl0_n_158, ZN => lbl0_d_position_1(0));
  lbl0_g18634 : AOI22D0BWP7T port map(A1 => lbl0_n_243, A2 => lbl0_n_125, B1 => lbl0_n_121, B2 => lbl0_n_117, ZN => lbl0_n_276);
  lbl0_g18635 : AOI21D0BWP7T port map(A1 => lbl0_n_175, A2 => lbl0_state(2), B => lbl0_n_254, ZN => lbl0_n_275);
  lbl0_g18636 : AOI32D0BWP7T port map(A1 => lbl0_n_121, A2 => lbl0_n_119, A3 => lbl0_n_85, B1 => lbl0_n_243, B2 => lbl0_n_109, ZN => lbl0_n_274);
  lbl0_g18637 : AOI211D0BWP7T port map(A1 => lbl0_n_217, A2 => lbl0_n_72, B => lbl0_n_221, C => lbl0_n_532, ZN => lbl0_n_273);
  lbl0_g18638 : OAI211D1BWP7T port map(A1 => lbl0_n_94, A2 => lbl0_n_103, B => lbl0_n_244, C => lbl0_n_122, ZN => lbl0_n_272);
  lbl0_g18639 : OAI31D0BWP7T port map(A1 => lbl0_state(2), A2 => lbl0_n_105, A3 => lbl0_n_172, B => lbl0_n_261, ZN => lbl0_n_281);
  lbl0_g18640 : MUX2ND0BWP7T port map(I0 => lbl0_n_53, I1 => lbl0_n_238, S => position_1(3), ZN => lbl0_n_280);
  lbl0_g18641 : IND3D0BWP7T port map(A1 => lbl0_n_439, B1 => lbl0_busy_count(6), B2 => lbl0_busy_count(5), ZN => lbl0_n_279);
  lbl0_g18642 : AOI21D0BWP7T port map(A1 => lbl0_n_141, A2 => lbl0_n_139, B => lbl0_n_267, ZN => lbl0_n_278);
  lbl0_g18643 : OAI21D0BWP7T port map(A1 => lbl0_n_532, A2 => lbl0_n_148, B => lbl0_n_266, ZN => lbl0_n_277);
  lbl0_g18645 : INVD1BWP7T port map(I => lbl0_n_266, ZN => lbl0_n_267);
  lbl0_g18646 : AOI221D0BWP7T port map(A1 => borders(0), A2 => lbl0_n_114, B1 => borders(1), B2 => lbl0_n_93, C => lbl0_n_225, ZN => lbl0_n_265);
  lbl0_g18647 : AN2D0BWP7T port map(A1 => lbl0_n_451, A2 => FE_PHN253_direction_between_3, Z => lbl0_d_next_direction_1(1));
  lbl0_g18648 : IND2D1BWP7T port map(A1 => lbl0_n_453, B1 => lbl0_n_248, ZN => lbl0_d_move_0);
  lbl0_g18649 : IND2D1BWP7T port map(A1 => lbl0_n_454, B1 => lbl0_n_248, ZN => lbl0_d_move_1);
  lbl0_g18650 : AN2D0BWP7T port map(A1 => lbl0_n_452, A2 => FE_PHN240_direction_between_0, Z => lbl0_d_next_direction_0(0));
  lbl0_g18651 : AN2D0BWP7T port map(A1 => lbl0_n_451, A2 => FE_PHN241_direction_between_2, Z => lbl0_d_next_direction_1(0));
  lbl0_g18652 : AN2D0BWP7T port map(A1 => lbl0_n_452, A2 => FE_PHN218_direction_between_1, Z => lbl0_d_next_direction_0(1));
  lbl0_g18653 : ND2D1BWP7T port map(A1 => lbl0_n_181, A2 => lbl0_n_226, ZN => lbl0_n_264);
  lbl0_g18654 : AOI221D0BWP7T port map(A1 => ramps(0), A2 => lbl0_n_91, B1 => ramps(1), B2 => lbl0_n_98, C => lbl0_n_227, ZN => lbl0_n_263);
  lbl0_g18655 : NR2D0BWP7T port map(A1 => lbl0_n_240, A2 => lbl0_n_52, ZN => lbl0_n_262);
  lbl0_g18656 : IND2D1BWP7T port map(A1 => lbl0_n_141, B1 => lbl0_n_450, ZN => lbl0_n_271);
  lbl0_g18657 : ND2D1BWP7T port map(A1 => lbl0_n_450, A2 => lbl0_n_148, ZN => lbl0_n_270);
  lbl0_g18658 : NR2D1BWP7T port map(A1 => lbl0_n_53, A2 => lbl0_n_238, ZN => lbl0_n_269);
  lbl0_g18659 : NR3D0BWP7T port map(A1 => lbl0_n_130, A2 => lbl0_n_66, A3 => FE_PHN262_lbl0_mem_com_state_3, ZN => lbl0_n_268);
  lbl0_g18660 : AOI211XD0BWP7T port map(A1 => lbl0_n_104, A2 => lbl0_n_79, B => lbl0_n_153, C => FE_PHN262_lbl0_mem_com_state_3, ZN => lbl0_n_266);
  lbl0_g18661 : INVD0BWP7T port map(I => lbl0_n_256, ZN => lbl0_n_255);
  lbl0_g18662 : OAI22D0BWP7T port map(A1 => lbl0_n_189, A2 => lbl0_move_1, B1 => lbl0_n_102, B2 => lbl0_n_94, ZN => lbl0_n_254);
  lbl0_g18663 : ND3D0BWP7T port map(A1 => lbl0_n_188, A2 => lbl0_n_149, A3 => lbl0_n_101, ZN => game_state(0));
  lbl0_g18664 : OAI221D0BWP7T port map(A1 => lbl0_n_174, A2 => lbl0_n_92, B1 => lbl0_n_116, B2 => lbl0_n_165, C => lbl0_next_direction_0(0), ZN => lbl0_n_253);
  lbl0_g18665 : MAOI22D0BWP7T port map(A1 => lbl0_n_185, A2 => lbl0_n_90, B1 => ramps(4), B2 => lbl0_n_90, ZN => lbl0_n_252);
  lbl0_g18666 : OAI21D0BWP7T port map(A1 => lbl0_n_208, A2 => FE_PHN207_lbl0_n_81, B => lbl0_n_158, ZN => lbl0_d_layer_1);
  lbl0_g18667 : AO21D0BWP7T port map(A1 => lbl0_n_104, A2 => lbl0_mem_com_state(1), B => lbl0_n_192, Z => write_enable);
  lbl0_g18668 : OAI21D0BWP7T port map(A1 => lbl0_n_207, A2 => FE_PHN210_lbl0_n_65, B => lbl0_n_158, ZN => lbl0_d_layer_0);
  lbl0_g18669 : AOI221D0BWP7T port map(A1 => ramps(2), A2 => lbl0_n_163, B1 => ramps(3), B2 => lbl0_n_115, C => lbl0_n_182, ZN => lbl0_n_251);
  lbl0_g18670 : AOI222D0BWP7T port map(A1 => lbl0_busy_count(2), A2 => lbl0_n_71, B1 => lbl0_n_129, B2 => lbl0_n_503, C1 => lbl0_n_112, C2 => lbl0_busy_count(1), ZN => lbl0_n_250);
  lbl0_g18671 : MOAI22D0BWP7T port map(A1 => lbl0_n_208, A2 => lbl0_n_137, B1 => lbl0_n_157, B2 => start_position_1(5), ZN => lbl0_d_position_1(5));
  lbl0_g18672 : OA33D0BWP7T port map(A1 => lbl0_n_59, A2 => lbl0_n_97, A3 => lbl0_n_172, B1 => lbl0_n_85, B2 => lbl0_state(3), B3 => lbl0_n_158, Z => lbl0_n_261);
  lbl0_g18673 : MOAI22D0BWP7T port map(A1 => lbl0_n_195, A2 => position_0(6), B1 => lbl0_n_195, B2 => position_0(6), ZN => lbl0_n_260);
  lbl0_g18674 : MOAI22D0BWP7T port map(A1 => lbl0_n_202, A2 => position_1(5), B1 => lbl0_n_202, B2 => position_1(5), ZN => lbl0_n_259);
  lbl0_g18675 : AO32D1BWP7T port map(A1 => lbl0_n_165, A2 => lbl0_n_115, A3 => position_0(3), B1 => lbl0_n_190, B2 => lbl0_n_83, Z => lbl0_n_258);
  lbl0_g18676 : AOI221D0BWP7T port map(A1 => lbl0_n_76, A2 => position_0(1), B1 => lbl0_n_178, B2 => lbl0_n_93, C => lbl0_n_184, ZN => lbl0_n_257);
  lbl0_g18677 : MOAI22D0BWP7T port map(A1 => lbl0_n_219, A2 => position_1(1), B1 => lbl0_n_219, B2 => position_1(1), ZN => lbl0_n_256);
  lbl0_g18678 : INVD0BWP7T port map(I => lbl0_n_244, ZN => lbl0_n_449);
  lbl0_g18679 : NR2XD0BWP7T port map(A1 => lbl0_n_123, A2 => lbl0_n_66, ZN => clear_memory);
  lbl0_g18680 : INR2D1BWP7T port map(A1 => direction_between(2), B1 => lbl0_n_209, ZN => lbl0_d_speed_select(0));
  lbl0_g18681 : NR4D0BWP7T port map(A1 => lbl0_n_97, A2 => lbl0_n_101, A3 => lbl0_state(3), A4 => start_between, ZN => lbl0_n_242);
  lbl0_g18682 : INR2D1BWP7T port map(A1 => lbl0_n_533, B1 => FE_PHN61_lbl0_booster_sync, ZN => lbl0_d_booster_sync);
  lbl0_g18683 : OR2D1BWP7T port map(A1 => lbl0_n_192, A2 => lbl0_mem_com_n_175, Z => go_to);
  lbl0_g18684 : INR2D1BWP7T port map(A1 => FE_PHN253_direction_between_3, B1 => lbl0_n_209, ZN => lbl0_d_speed_select(1));
  lbl0_g18685 : INR2D1BWP7T port map(A1 => lbl0_n_136, B1 => lbl0_n_207, ZN => lbl0_n_442);
  lbl0_g18686 : INR2D1BWP7T port map(A1 => FE_PHN240_direction_between_0, B1 => lbl0_n_209, ZN => lbl0_d_map_select(0));
  lbl0_g18687 : NR2D1BWP7T port map(A1 => lbl0_n_207, A2 => lbl0_n_135, ZN => lbl0_n_440);
  lbl0_g18688 : INR2D1BWP7T port map(A1 => FE_PHN218_direction_between_1, B1 => lbl0_n_209, ZN => lbl0_d_map_select(1));
  lbl0_g18689 : OR2D1BWP7T port map(A1 => lbl0_n_533, A2 => lbl0_n_157, Z => lbl0_n_456);
  lbl0_g18690 : NR2D0BWP7T port map(A1 => lbl0_n_218, A2 => lbl0_n_72, ZN => lbl0_n_249);
  lbl0_g18691 : ND2D1BWP7T port map(A1 => lbl0_n_533, A2 => FE_PHN61_lbl0_booster_sync, ZN => lbl0_n_248);
  lbl0_g18692 : ND2D0BWP7T port map(A1 => lbl0_n_535, A2 => start_between, ZN => lbl0_n_247);
  lbl0_g18693 : INR2D0BWP7T port map(A1 => lbl0_n_177, B1 => lbl0_n_220, ZN => lbl0_n_246);
  lbl0_g18695 : IND2D0BWP7T port map(A1 => lbl0_n_189, B1 => lbl0_move_0, ZN => lbl0_n_245);
  lbl0_g18696 : IND2D1BWP7T port map(A1 => lbl0_n_532, B1 => lbl0_n_139, ZN => lbl0_n_455);
  lbl0_g18698 : AN2D1BWP7T port map(A1 => lbl0_n_533, A2 => lbl0_n_201, Z => lbl0_n_451);
  lbl0_g18699 : AN2D1BWP7T port map(A1 => lbl0_n_533, A2 => lbl0_n_200, Z => lbl0_n_452);
  lbl0_g18700 : INR2XD0BWP7T port map(A1 => lbl0_n_191, B1 => lbl0_n_536, ZN => lbl0_n_244);
  lbl0_g18701 : OR2D1BWP7T port map(A1 => lbl0_n_446, A2 => lbl0_n_192, Z => lbl0_n_450);
  lbl0_g18702 : NR2D0BWP7T port map(A1 => lbl0_n_220, A2 => lbl0_n_177, ZN => lbl0_n_243);
  lbl0_g18703 : OR2D1BWP7T port map(A1 => lbl0_n_436, A2 => lbl0_n_2, Z => lbl0_n_439);
  lbl0_g18704 : INVD0BWP7T port map(I => lbl0_n_237, ZN => lbl0_n_236);
  lbl0_g18705 : OAI21D0BWP7T port map(A1 => lbl0_n_160, A2 => lbl0_n_76, B => lbl0_n_210, ZN => lbl0_d_direction_0(0));
  lbl0_g18706 : OAI221D0BWP7T port map(A1 => lbl0_n_92, A2 => lbl0_n_107, B1 => lbl0_n_116, B2 => lbl0_n_120, C => lbl0_next_direction_0(0), ZN => lbl0_n_235);
  lbl0_g18707 : AO211D0BWP7T port map(A1 => lbl0_n_98, A2 => position_1(1), B => lbl0_n_219, C => lbl0_n_156, Z => lbl0_n_234);
  lbl0_g18708 : MOAI22D0BWP7T port map(A1 => lbl0_n_136, A2 => lbl0_n_78, B1 => lbl0_n_136, B2 => lbl0_n_78, ZN => lbl0_n_233);
  lbl0_g18709 : ND3D0BWP7T port map(A1 => lbl0_n_175, A2 => lbl0_n_154, A3 => lbl0_n_94, ZN => game_state(2));
  lbl0_g18710 : OAI21D0BWP7T port map(A1 => lbl0_n_160, A2 => lbl0_n_55, B => lbl0_n_210, ZN => lbl0_d_direction_1(0));
  lbl0_g18711 : OA21D0BWP7T port map(A1 => lbl0_n_160, A2 => lbl0_n_151, B => lbl0_n_457, Z => lbl0_e_position_1);
  lbl0_g18712 : OA21D0BWP7T port map(A1 => lbl0_n_160, A2 => lbl0_n_144, B => lbl0_n_457, Z => lbl0_e_position_0);
  lbl0_g18713 : IOA21D1BWP7T port map(A1 => lbl0_n_159, A2 => FE_PHN196_lbl0_next_direction_0_1, B => lbl0_n_158, ZN => lbl0_d_direction_0(1));
  lbl0_g18715 : OAI22D0BWP7T port map(A1 => ramps(6), A2 => lbl0_n_162, B1 => ramps(7), B2 => lbl0_n_116, ZN => lbl0_n_232);
  lbl0_g18716 : AOI21D0BWP7T port map(A1 => lbl0_n_56, A2 => lbl0_move_0, B => lbl0_n_214, ZN => lbl0_n_231);
  lbl0_g18717 : AO21D0BWP7T port map(A1 => lbl0_n_165, A2 => lbl0_n_115, B => lbl0_n_190, Z => lbl0_n_230);
  lbl0_g18718 : IND3D1BWP7T port map(A1 => lbl0_n_166, B1 => lbl0_n_105, B2 => lbl0_n_149, ZN => game_state(1));
  lbl0_g18719 : AOI222D0BWP7T port map(A1 => borders(4), A2 => lbl0_n_91, B1 => borders(7), B2 => lbl0_n_96, C1 => borders(5), C2 => lbl0_n_98, ZN => lbl0_n_229);
  lbl0_g18720 : AOI222D0BWP7T port map(A1 => borders(0), A2 => lbl0_n_91, B1 => borders(3), B2 => lbl0_n_96, C1 => borders(1), C2 => lbl0_n_98, ZN => lbl0_n_228);
  lbl0_g18721 : AO32D1BWP7T port map(A1 => ramps(2), A2 => lbl0_n_90, A3 => lbl0_n_55, B1 => ramps(3), B2 => lbl0_n_96, Z => lbl0_n_227);
  lbl0_g18722 : AOI22D0BWP7T port map(A1 => borders(6), A2 => lbl0_n_163, B1 => borders(7), B2 => lbl0_n_115, ZN => lbl0_n_226);
  lbl0_g18723 : AO22D0BWP7T port map(A1 => borders(2), A2 => lbl0_n_163, B1 => lbl0_n_115, B2 => borders(3), Z => lbl0_n_225);
  lbl0_g18724 : OAI222D0BWP7T port map(A1 => lbl0_n_87, A2 => lbl0_next_direction_1(1), B1 => direction_1(0), B2 => lbl0_next_direction_1(0), C1 => direction_1(1), C2 => lbl0_n_63, ZN => lbl0_n_241);
  lbl0_g18725 : IND3D1BWP7T port map(A1 => lbl0_n_191, B1 => lbl0_n_152, B2 => lbl0_n_146, ZN => lbl0_n_240);
  lbl0_g18726 : OAI222D0BWP7T port map(A1 => lbl0_n_86, A2 => lbl0_next_direction_0(1), B1 => direction_0(0), B2 => lbl0_next_direction_0(0), C1 => direction_0(1), C2 => lbl0_n_62, ZN => lbl0_n_239);
  lbl0_g18727 : AN3D1BWP7T port map(A1 => lbl0_n_171, A2 => position_1(1), A3 => position_1(2), Z => lbl0_n_238);
  lbl0_g18729 : AOI211XD0BWP7T port map(A1 => lbl0_n_55, A2 => position_1(0), B => lbl0_n_169, C => lbl0_n_155, ZN => lbl0_n_237);
  lbl0_g18730 : CKND1BWP7T port map(I => lbl0_n_217, ZN => lbl0_n_218);
  lbl0_g18731 : INVD0BWP7T port map(I => lbl0_n_213, ZN => lbl0_n_212);
  lbl0_g18732 : INVD0BWP7T port map(I => lbl0_n_211, ZN => lbl0_n_210);
  lbl0_g18733 : INVD1BWP7T port map(I => lbl0_n_535, ZN => lbl0_n_209);
  lbl0_g18734 : INVD0BWP7T port map(I => lbl0_n_207, ZN => lbl0_n_206);
  lbl0_g18736 : NR2D1BWP7T port map(A1 => lbl0_n_164, A2 => lbl0_n_56, ZN => lbl0_n_531);
  lbl0_g18737 : NR2D1BWP7T port map(A1 => lbl0_n_160, A2 => FE_PHN167_lbl0_n_63, ZN => lbl0_d_direction_1(1));
  lbl0_g18738 : NR2XD0BWP7T port map(A1 => lbl0_n_173, A2 => lbl0_mem_com_state(1), ZN => lbl0_mem_com_n_166);
  lbl0_g18739 : OR2D1BWP7T port map(A1 => lbl0_n_134, A2 => lbl0_n_91, Z => lbl0_n_205);
  lbl0_g18740 : ND2D1BWP7T port map(A1 => lbl0_n_138, A2 => FE_PHN163_lbl0_border_0, ZN => lbl0_n_224);
  lbl0_g18741 : IND2D0BWP7T port map(A1 => lbl0_n_139, B1 => lbl0_n_59, ZN => lbl0_n_223);
  lbl0_g18742 : ND2D1BWP7T port map(A1 => lbl0_n_138, A2 => FE_PHN340_lbl0_border_1, ZN => lbl0_n_222);
  lbl0_g18743 : NR2XD0BWP7T port map(A1 => lbl0_n_173, A2 => lbl0_n_79, ZN => lbl0_n_446);
  lbl0_g18744 : NR2D0BWP7T port map(A1 => lbl0_n_167, A2 => lbl0_n_97, ZN => lbl0_n_221);
  lbl0_g18745 : IND2D0BWP7T port map(A1 => lbl0_n_97, B1 => lbl0_n_176, ZN => lbl0_n_220);
  lbl0_g18746 : NR2D1BWP7T port map(A1 => lbl0_n_169, A2 => lbl0_n_171, ZN => lbl0_n_219);
  lbl0_g18747 : NR2D0BWP7T port map(A1 => lbl0_n_142, A2 => lbl0_state(4), ZN => lbl0_n_217);
  lbl0_g18748 : AN2D1BWP7T port map(A1 => lbl0_n_161, A2 => lbl0_n_119, Z => lbl0_n_536);
  lbl0_g18749 : ND2D0BWP7T port map(A1 => lbl0_n_176, A2 => lbl0_state(2), ZN => lbl0_n_216);
  lbl0_g18750 : ND2D1BWP7T port map(A1 => lbl0_n_160, A2 => lbl0_n_158, ZN => lbl0_n_457);
  lbl0_g18751 : ND2D1BWP7T port map(A1 => lbl0_n_157, A2 => start_position_0(2), ZN => lbl0_n_215);
  lbl0_g18752 : ND2D0BWP7T port map(A1 => lbl0_n_166, A2 => lbl0_state(3), ZN => lbl0_n_214);
  lbl0_g18753 : IND2D1BWP7T port map(A1 => lbl0_n_94, B1 => lbl0_n_161, ZN => lbl0_n_213);
  lbl0_g18754 : AN2D1BWP7T port map(A1 => lbl0_n_161, A2 => lbl0_n_117, Z => lbl0_n_532);
  lbl0_g18755 : NR2D1BWP7T port map(A1 => lbl0_n_158, A2 => start_position_0(2), ZN => lbl0_n_211);
  lbl0_g18756 : INR2D1BWP7T port map(A1 => lbl0_n_161, B1 => lbl0_n_97, ZN => lbl0_n_535);
  lbl0_g18757 : NR2XD0BWP7T port map(A1 => lbl0_n_168, A2 => lbl0_n_118, ZN => lbl0_n_533);
  lbl0_g18758 : ND2D1BWP7T port map(A1 => lbl0_n_159, A2 => lbl0_n_151, ZN => lbl0_n_208);
  lbl0_g18759 : ND2D1BWP7T port map(A1 => lbl0_n_159, A2 => lbl0_n_144, ZN => lbl0_n_207);
  lbl0_g18762 : INVD0BWP7T port map(I => lbl0_n_198, ZN => lbl0_n_199);
  lbl0_g18763 : INVD0BWP7T port map(I => lbl0_n_196, ZN => lbl0_n_197);
  lbl0_g18764 : MAOI22D0BWP7T port map(A1 => lbl0_n_111, A2 => lbl0_state(2), B1 => lbl0_n_111, B2 => lbl0_state(2), ZN => lbl0_n_188);
  lbl0_g18765 : NR4D0BWP7T port map(A1 => read_memory_in(3), A2 => read_memory_in(2), A3 => read_memory_in(1), A4 => read_memory_in(0), ZN => lbl0_n_187);
  lbl0_g18766 : AN3D0BWP7T port map(A1 => lbl0_n_120, A2 => lbl0_n_115, A3 => lbl0_n_80, Z => lbl0_n_186);
  lbl0_g18767 : NR3D0BWP7T port map(A1 => ramps(6), A2 => lbl0_n_96, A3 => lbl0_n_98, ZN => lbl0_n_185);
  lbl0_g18768 : NR2D0BWP7T port map(A1 => lbl0_n_178, A2 => lbl0_n_116, ZN => lbl0_n_184);
  lbl0_g18769 : OAI22D0BWP7T port map(A1 => ramps(4), A2 => lbl0_n_113, B1 => ramps(5), B2 => lbl0_n_92, ZN => lbl0_n_183);
  lbl0_g18770 : AO22D0BWP7T port map(A1 => ramps(0), A2 => lbl0_n_114, B1 => lbl0_n_93, B2 => ramps(1), Z => lbl0_n_182);
  lbl0_g18771 : AOI22D0BWP7T port map(A1 => borders(4), A2 => lbl0_n_114, B1 => borders(5), B2 => lbl0_n_93, ZN => lbl0_n_181);
  lbl0_g18772 : NR4D0BWP7T port map(A1 => read_memory_in(7), A2 => read_memory_in(6), A3 => read_memory_in(5), A4 => read_memory_in(4), ZN => lbl0_n_180);
  lbl0_g18773 : MOAI22D0BWP7T port map(A1 => lbl0_n_90, A2 => position_1(9), B1 => lbl0_n_90, B2 => position_1(9), ZN => lbl0_n_204);
  lbl0_g18774 : MOAI22D0BWP7T port map(A1 => lbl0_n_90, A2 => position_1(7), B1 => lbl0_n_90, B2 => position_1(7), ZN => lbl0_n_203);
  lbl0_g18775 : MAOI22D0BWP7T port map(A1 => lbl0_n_90, A2 => position_1(6), B1 => lbl0_n_90, B2 => position_1(6), ZN => lbl0_n_202);
  lbl0_g18777 : ND2D1BWP7T port map(A1 => lbl0_n_145, A2 => lbl0_n_143, ZN => lbl0_n_201);
  lbl0_g18778 : IND2D1BWP7T port map(A1 => lbl0_n_146, B1 => lbl0_n_152, ZN => lbl0_n_200);
  lbl0_g18779 : IND3D1BWP7T port map(A1 => lbl0_n_437, B1 => lbl0_busy_count(2), B2 => lbl0_busy_count(3), ZN => lbl0_n_436);
  lbl0_g18780 : MOAI22D0BWP7T port map(A1 => lbl0_n_127, A2 => lbl0_n_110, B1 => lbl0_n_127, B2 => lbl0_n_110, ZN => lbl0_n_198);
  lbl0_g18781 : MOAI22D0BWP7T port map(A1 => lbl0_n_108, A2 => lbl0_n_124, B1 => lbl0_n_108, B2 => lbl0_n_124, ZN => lbl0_n_196);
  lbl0_g18782 : MAOI22D0BWP7T port map(A1 => lbl0_n_113, A2 => position_0(5), B1 => lbl0_n_113, B2 => position_0(5), ZN => lbl0_n_195);
  lbl0_g18783 : MAOI222D1BWP7T port map(A => lbl0_n_114, B => position_0(6), C => position_0(5), ZN => lbl0_n_194);
  lbl0_g18784 : MAOI222D1BWP7T port map(A => lbl0_n_91, B => position_1(6), C => position_1(5), ZN => lbl0_n_193);
  lbl0_g18785 : NR4D0BWP7T port map(A1 => lbl0_n_67, A2 => lbl0_mem_com_state(2), A3 => lbl0_mem_com_state(1), A4 => FE_PHN262_lbl0_mem_com_state_3, ZN => lbl0_n_192);
  lbl0_g18786 : OR2D1BWP7T port map(A1 => lbl0_n_168, A2 => lbl0_n_94, Z => lbl0_n_191);
  lbl0_g18787 : AN2D1BWP7T port map(A1 => lbl0_n_174, A2 => lbl0_n_93, Z => lbl0_n_190);
  lbl0_g18788 : OR2D0BWP7T port map(A1 => lbl0_n_168, A2 => lbl0_n_97, Z => lbl0_n_189);
  lbl0_g18789 : CKND1BWP7T port map(I => lbl0_n_170, ZN => lbl0_n_171);
  lbl0_g18791 : INVD0BWP7T port map(I => lbl0_n_163, ZN => lbl0_n_162);
  lbl0_g18792 : INVD1BWP7T port map(I => lbl0_n_160, ZN => lbl0_n_159);
  lbl0_g18793 : INVD1BWP7T port map(I => lbl0_n_158, ZN => lbl0_n_157);
  lbl0_g18794 : NR2D0BWP7T port map(A1 => lbl0_n_95, A2 => position_1(1), ZN => lbl0_n_156);
  lbl0_g18795 : NR2D1BWP7T port map(A1 => lbl0_n_95, A2 => position_1(0), ZN => lbl0_n_155);
  lbl0_g18796 : ND2D1BWP7T port map(A1 => lbl0_n_97, A2 => lbl0_n_122, ZN => lbl0_n_154);
  lbl0_g18797 : NR2D1BWP7T port map(A1 => lbl0_n_104, A2 => lbl0_n_79, ZN => lbl0_n_153);
  lbl0_g18798 : IND2D0BWP7T port map(A1 => lbl0_n_105, B1 => lbl0_n_121, ZN => lbl0_n_179);
  lbl0_g18799 : OR2D0BWP7T port map(A1 => lbl0_n_120, A2 => lbl0_n_107, Z => lbl0_n_178);
  lbl0_g18800 : NR2D0BWP7T port map(A1 => lbl0_n_109, A2 => lbl0_n_125, ZN => lbl0_n_177);
  lbl0_g18801 : INR2D0BWP7T port map(A1 => lbl0_n_100, B1 => lbl0_state(4), ZN => lbl0_n_176);
  lbl0_g18802 : CKAN2D1BWP7T port map(A1 => lbl0_n_102, A2 => lbl0_n_58, Z => lbl0_n_175);
  lbl0_g18803 : CKAN2D1BWP7T port map(A1 => lbl0_n_107, A2 => lbl0_n_80, Z => lbl0_n_174);
  lbl0_g18804 : IND2D1BWP7T port map(A1 => FE_PHN262_lbl0_mem_com_state_3, B1 => lbl0_n_104, ZN => lbl0_n_173);
  lbl0_g18805 : NR2XD0BWP7T port map(A1 => lbl0_n_126, A2 => lbl0_mem_com_state(1), ZN => lbl0_mem_com_n_175);
  lbl0_g18806 : IND2D0BWP7T port map(A1 => lbl0_n_106, B1 => lbl0_n_85, ZN => lbl0_n_172);
  lbl0_g18807 : ND2D1BWP7T port map(A1 => lbl0_n_96, A2 => position_1(0), ZN => lbl0_n_170);
  lbl0_g18808 : NR2XD0BWP7T port map(A1 => lbl0_n_99, A2 => position_1(0), ZN => lbl0_n_169);
  lbl0_g18809 : OR2D1BWP7T port map(A1 => lbl0_n_102, A2 => lbl0_state(3), Z => lbl0_n_168);
  lbl0_g18810 : IND2D0BWP7T port map(A1 => lbl0_n_102, B1 => lbl0_state(3), ZN => lbl0_n_167);
  lbl0_g18811 : NR2D1BWP7T port map(A1 => lbl0_n_118, A2 => lbl0_state(4), ZN => lbl0_n_166);
  lbl0_g18812 : CKAN2D1BWP7T port map(A1 => lbl0_n_120, A2 => position_0(2), Z => lbl0_n_165);
  lbl0_g18813 : OR2D1BWP7T port map(A1 => lbl0_n_105, A2 => lbl0_n_5, Z => lbl0_n_164);
  lbl0_g18814 : NR2D1BWP7T port map(A1 => lbl0_n_114, A2 => lbl0_next_direction_0(0), ZN => lbl0_n_163);
  lbl0_g18815 : NR2D1BWP7T port map(A1 => lbl0_n_106, A2 => lbl0_state(4), ZN => lbl0_n_161);
  lbl0_g18816 : ND2D1BWP7T port map(A1 => lbl0_n_100, A2 => lbl0_n_117, ZN => lbl0_n_160);
  lbl0_g18817 : OR2D1BWP7T port map(A1 => lbl0_n_122, A2 => lbl0_n_118, Z => lbl0_n_158);
  lbl0_g18819 : AOI22D0BWP7T port map(A1 => borders(2), A2 => FE_DBTN22_position_1_10, B1 => borders(6), B2 => position_1(10), ZN => lbl0_n_134);
  lbl0_g18820 : AOI22D0BWP7T port map(A1 => lbl0_n_65, A2 => position_1(10), B1 => FE_DBTN22_position_1_10, B2 => lbl0_next_layer_0, ZN => lbl0_n_133);
  lbl0_g18821 : MAOI22D0BWP7T port map(A1 => lbl0_n_81, A2 => position_0(10), B1 => lbl0_n_81, B2 => position_0(10), ZN => lbl0_n_132);
  lbl0_g18822 : AOI22D0BWP7T port map(A1 => lbl0_n_81, A2 => lbl0_n_65, B1 => lbl0_next_layer_0, B2 => lbl0_next_layer_1, ZN => lbl0_n_131);
  lbl0_g18823 : OAI21D0BWP7T port map(A1 => lbl0_mem_com_state(0), A2 => lbl0_mem_com_state(1), B => lbl0_n_123, ZN => lbl0_n_130);
  lbl0_g18824 : IOA21D0BWP7T port map(A1 => FE_PHN258_lbl0_busy_count_0, A2 => lbl0_busy_count(2), B => lbl0_n_502, ZN => lbl0_n_129);
  lbl0_g18825 : MOAI22D0BWP7T port map(A1 => direction_0(0), A2 => FE_PHN240_direction_between_0, B1 => direction_0(0), B2 => FE_PHN240_direction_between_0, ZN => lbl0_n_152);
  lbl0_g18826 : AOI21D0BWP7T port map(A1 => lbl0_n_89, A2 => player_state_1(0), B => lbl0_n_72, ZN => lbl0_n_151);
  lbl0_g18827 : MOAI22D0BWP7T port map(A1 => lbl0_n_55, A2 => direction_1(0), B1 => lbl0_n_55, B2 => direction_1(0), ZN => lbl0_n_150);
  lbl0_g18828 : AOI21D0BWP7T port map(A1 => lbl0_n_56, A2 => lbl0_state(1), B => lbl0_state(3), ZN => lbl0_n_149);
  lbl0_g18829 : NR2D1BWP7T port map(A1 => lbl0_n_101, A2 => lbl0_n_118, ZN => lbl0_n_530);
  lbl0_g18830 : INR2D1BWP7T port map(A1 => lbl0_n_100, B1 => lbl0_n_94, ZN => lbl0_n_148);
  lbl0_g18831 : MOAI22D0BWP7T port map(A1 => lbl0_n_76, A2 => direction_0(0), B1 => lbl0_n_76, B2 => direction_0(0), ZN => lbl0_n_147);
  lbl0_g18832 : MOAI22D0BWP7T port map(A1 => direction_0(1), A2 => direction_between(1), B1 => direction_0(1), B2 => direction_between(1), ZN => lbl0_n_146);
  lbl0_g18833 : MAOI22D0BWP7T port map(A1 => direction_1(1), A2 => FE_PHN253_direction_between_3, B1 => direction_1(1), B2 => FE_PHN253_direction_between_3, ZN => lbl0_n_145);
  lbl0_g18834 : OA21D0BWP7T port map(A1 => lbl0_n_88, A2 => player_state_0(1), B => lbl0_move_0, Z => lbl0_n_144);
  lbl0_g18835 : MOAI22D0BWP7T port map(A1 => direction_1(0), A2 => direction_between(2), B1 => direction_1(0), B2 => direction_between(2), ZN => lbl0_n_143);
  lbl0_g18836 : ND2D1BWP7T port map(A1 => lbl0_n_100, A2 => lbl0_n_119, ZN => lbl0_n_142);
  lbl0_g18837 : OR2D1BWP7T port map(A1 => lbl0_n_103, A2 => lbl0_n_118, Z => lbl0_n_141);
  lbl0_g18838 : OR2D1BWP7T port map(A1 => lbl0_n_103, A2 => lbl0_n_97, Z => lbl0_n_140);
  lbl0_g18839 : IND2D1BWP7T port map(A1 => lbl0_n_103, B1 => lbl0_n_119, ZN => lbl0_n_139);
  lbl0_g18840 : INR2XD0BWP7T port map(A1 => lbl0_n_119, B1 => lbl0_n_101, ZN => lbl0_n_138);
  lbl0_g18841 : AOI22D0BWP7T port map(A1 => lbl0_n_55, A2 => lbl0_n_78, B1 => lbl0_next_direction_1(0), B2 => position_1(5), ZN => lbl0_n_137);
  lbl0_g18842 : MOAI22D0BWP7T port map(A1 => lbl0_next_direction_0(0), A2 => position_0(5), B1 => lbl0_next_direction_0(0), B2 => position_0(5), ZN => lbl0_n_136);
  lbl0_g18843 : AOI22D0BWP7T port map(A1 => lbl0_n_82, A2 => lbl0_next_direction_0(0), B1 => lbl0_n_76, B2 => position_0(0), ZN => lbl0_n_135);
  lbl0_g18845 : INVD0BWP7T port map(I => lbl0_n_118, ZN => lbl0_n_117);
  lbl0_g18846 : INVD1BWP7T port map(I => lbl0_n_116, ZN => lbl0_n_115);
  lbl0_g18847 : INVD1BWP7T port map(I => lbl0_n_114, ZN => lbl0_n_113);
  lbl0_g18848 : CKAN2D1BWP7T port map(A1 => lbl0_busy_count(4), A2 => lbl0_busy_count(5), Z => lbl0_n_438);
  lbl0_g18849 : ND2D0BWP7T port map(A1 => lbl0_state(0), A2 => lbl0_state(1), ZN => lbl0_n_461);
  lbl0_g18850 : ND2D0BWP7T port map(A1 => lbl0_n_4, A2 => lbl0_n_502, ZN => lbl0_n_112);
  lbl0_g18851 : CKND2D1BWP7T port map(A1 => lbl0_mem_com_state(0), A2 => FE_PHN262_lbl0_mem_com_state_3, ZN => lbl0_n_128);
  lbl0_g18852 : NR2D1BWP7T port map(A1 => lbl0_next_direction_0(0), A2 => direction_0(1), ZN => lbl0_n_127);
  lbl0_g18853 : ND2D1BWP7T port map(A1 => lbl0_n_67, A2 => lbl0_mem_com_state(2), ZN => lbl0_n_126);
  lbl0_g18854 : ND2D0BWP7T port map(A1 => player_state_0(0), A2 => player_state_0(1), ZN => lbl0_n_125);
  lbl0_g18855 : IND2D1BWP7T port map(A1 => direction_1(0), B1 => lbl0_next_direction_1(1), ZN => lbl0_n_124);
  lbl0_g18856 : ND2D1BWP7T port map(A1 => lbl0_mem_com_state(1), A2 => lbl0_mem_com_state(0), ZN => lbl0_n_123);
  lbl0_g18857 : CKND2D1BWP7T port map(A1 => FE_PHN258_lbl0_busy_count_0, A2 => lbl0_busy_count(1), ZN => lbl0_n_437);
  lbl0_g18858 : ND2D1BWP7T port map(A1 => lbl0_state(4), A2 => lbl0_state(0), ZN => lbl0_n_122);
  lbl0_g18859 : NR2D0BWP7T port map(A1 => lbl0_state(0), A2 => lbl0_state(3), ZN => lbl0_n_121);
  lbl0_g18860 : NR2XD0BWP7T port map(A1 => lbl0_n_82, A2 => lbl0_n_84, ZN => lbl0_n_120);
  lbl0_g18861 : NR2D1BWP7T port map(A1 => lbl0_state(2), A2 => lbl0_state(1), ZN => lbl0_n_119);
  lbl0_g18862 : ND2D1BWP7T port map(A1 => lbl0_state(1), A2 => lbl0_state(2), ZN => lbl0_n_118);
  lbl0_g18863 : CKND2D1BWP7T port map(A1 => lbl0_next_direction_0(1), A2 => lbl0_next_direction_0(0), ZN => lbl0_n_116);
  lbl0_g18864 : NR2XD0BWP7T port map(A1 => lbl0_next_direction_0(0), A2 => lbl0_next_direction_0(1), ZN => lbl0_n_114);
  lbl0_g18865 : INVD1BWP7T port map(I => lbl0_n_99, ZN => lbl0_n_98);
  lbl0_g18866 : INVD0BWP7T port map(I => lbl0_n_96, ZN => lbl0_n_95);
  lbl0_g18867 : INVD0BWP7T port map(I => lbl0_n_93, ZN => lbl0_n_92);
  lbl0_g18868 : INVD1BWP7T port map(I => lbl0_n_91, ZN => lbl0_n_90);
  lbl0_g18869 : ND2D1BWP7T port map(A1 => lbl0_state(1), A2 => lbl0_state(4), ZN => lbl0_n_111);
  lbl0_g18870 : IND2D1BWP7T port map(A1 => direction_0(0), B1 => lbl0_next_direction_0(1), ZN => lbl0_n_110);
  lbl0_g18871 : ND2D0BWP7T port map(A1 => player_state_1(0), A2 => player_state_1(1), ZN => lbl0_n_109);
  lbl0_g18872 : NR2D1BWP7T port map(A1 => lbl0_next_direction_1(0), A2 => direction_1(1), ZN => lbl0_n_108);
  lbl0_g18873 : NR2XD0BWP7T port map(A1 => position_0(1), A2 => position_0(0), ZN => lbl0_n_107);
  lbl0_g18874 : CKND2D1BWP7T port map(A1 => lbl0_n_58, A2 => lbl0_state(0), ZN => lbl0_n_106);
  lbl0_g18875 : CKND2D1BWP7T port map(A1 => lbl0_n_60, A2 => lbl0_state(4), ZN => lbl0_n_105);
  lbl0_g18876 : NR2XD0BWP7T port map(A1 => lbl0_mem_com_state(2), A2 => lbl0_mem_com_state(0), ZN => lbl0_n_104);
  lbl0_g18877 : ND2D1BWP7T port map(A1 => lbl0_n_56, A2 => lbl0_state(3), ZN => lbl0_n_103);
  lbl0_g18878 : CKND2D1BWP7T port map(A1 => lbl0_n_59, A2 => lbl0_n_56, ZN => lbl0_n_102);
  lbl0_g18879 : CKND2D1BWP7T port map(A1 => lbl0_n_56, A2 => lbl0_state(4), ZN => lbl0_n_101);
  lbl0_g18880 : NR2D1BWP7T port map(A1 => lbl0_n_58, A2 => lbl0_n_56, ZN => lbl0_n_100);
  lbl0_g18881 : ND2D1BWP7T port map(A1 => lbl0_n_63, A2 => lbl0_next_direction_1(0), ZN => lbl0_n_99);
  lbl0_g18882 : ND2D1BWP7T port map(A1 => lbl0_n_5, A2 => lbl0_state(1), ZN => lbl0_n_97);
  lbl0_g18883 : NR2XD0BWP7T port map(A1 => lbl0_n_55, A2 => lbl0_n_63, ZN => lbl0_n_96);
  lbl0_g18884 : CKND2D1BWP7T port map(A1 => lbl0_n_60, A2 => lbl0_state(2), ZN => lbl0_n_94);
  lbl0_g18885 : NR2D1BWP7T port map(A1 => lbl0_n_76, A2 => lbl0_next_direction_0(1), ZN => lbl0_n_93);
  lbl0_g18886 : NR2XD0BWP7T port map(A1 => lbl0_next_direction_1(0), A2 => lbl0_next_direction_1(1), ZN => lbl0_n_91);
  lbl0_g18887 : INVD0BWP7T port map(I => player_state_1(1), ZN => lbl0_n_89);
  lbl0_g18888 : CKND1BWP7T port map(I => player_state_0(0), ZN => lbl0_n_88);
  lbl0_g18889 : INVD0BWP7T port map(I => direction_1(1), ZN => lbl0_n_87);
  lbl0_g18890 : INVD0BWP7T port map(I => direction_0(1), ZN => lbl0_n_86);
  lbl0_g18891 : INVD0BWP7T port map(I => start_between, ZN => lbl0_n_85);
  lbl0_g18892 : INVD1BWP7T port map(I => position_0(1), ZN => lbl0_n_84);
  lbl0_g18893 : INVD1BWP7T port map(I => position_0(3), ZN => lbl0_n_83);
  lbl0_g18894 : INVD1BWP7T port map(I => position_0(0), ZN => lbl0_n_82);
  lbl0_g18895 : INVD1BWP7T port map(I => lbl0_next_layer_1, ZN => lbl0_n_81);
  lbl0_g18896 : INVD0BWP7T port map(I => position_0(2), ZN => lbl0_n_80);
  lbl0_g18899 : INVD0BWP7T port map(I => position_1(5), ZN => lbl0_n_78);
  lbl0_g18901 : INVD1BWP7T port map(I => lbl0_next_direction_0(0), ZN => lbl0_n_76);
  lbl0_g18902 : INVD0BWP7T port map(I => lbl0_read_data_reg(7), ZN => lbl0_n_75);
  lbl0_g18903 : INVD0BWP7T port map(I => lbl0_read_data_reg(5), ZN => lbl0_n_74);
  lbl0_g18904 : INVD0BWP7T port map(I => lbl0_read_data_reg(4), ZN => lbl0_n_73);
  lbl0_g18905 : INVD1BWP7T port map(I => lbl0_move_1, ZN => lbl0_n_72);
  lbl0_g18906 : INVD0BWP7T port map(I => lbl0_n_502, ZN => lbl0_n_71);
  lbl0_g18909 : INVD1BWP7T port map(I => position_0(4), ZN => lbl0_n_68);
  lbl0_g18912 : INVD1BWP7T port map(I => lbl0_next_layer_0, ZN => lbl0_n_65);
  lbl0_g18913 : INVD1BWP7T port map(I => position_1(8), ZN => lbl0_n_64);
  lbl0_g18914 : INVD1BWP7T port map(I => lbl0_next_direction_1(1), ZN => lbl0_n_63);
  lbl0_g18915 : INVD0BWP7T port map(I => lbl0_next_direction_0(1), ZN => lbl0_n_62);
  lbl0_g18916 : INVD1BWP7T port map(I => position_0(7), ZN => lbl0_n_61);
  lbl0_g18922 : INVD1BWP7T port map(I => lbl0_next_direction_1(0), ZN => lbl0_n_55);
  lbl0_g2 : IND2D1BWP7T port map(A1 => lbl0_n_270, B1 => position_0(10), ZN => lbl0_n_54);
  lbl0_g18923 : INR2D1BWP7T port map(A1 => lbl0_n_533, B1 => lbl0_n_201, ZN => lbl0_n_454);
  lbl0_g18924 : INR2D1BWP7T port map(A1 => lbl0_n_533, B1 => lbl0_n_200, ZN => lbl0_n_453);
  lbl0_g18925 : INR3D0BWP7T port map(A1 => lbl0_n_169, B1 => position_1(1), B2 => position_1(2), ZN => lbl0_n_53);
  lbl0_g18926 : IND2D1BWP7T port map(A1 => lbl0_n_145, B1 => lbl0_n_143, ZN => lbl0_n_52);
  lbl0_g18927 : INR3D0BWP7T port map(A1 => position_1(1), B1 => lbl0_n_170, B2 => position_1(2), ZN => lbl0_n_51);
  lbl0_g8596 : ND4D0BWP7T port map(A1 => lbl0_n_542, A2 => lbl0_n_49, A3 => lbl0_n_22, A4 => FE_PHN309_lbl0_n_539, ZN => lbl0_n_50);
  lbl0_g8601 : MAOI22D0BWP7T port map(A1 => memory_ready, A2 => lbl0_n_41, B1 => lbl0_n_9, B2 => lbl0_n_28, ZN => lbl0_n_49);
  lbl0_mem_com_state_reg_3 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN311_lbl0_n_47, Q => lbl0_mem_com_state(3));
  lbl0_g8605 : ND2D1BWP7T port map(A1 => lbl0_n_40, A2 => lbl0_n_22, ZN => lbl0_n_48);
  lbl0_counter_busy_counter_state_reg_0 : DFKCNQD1BWP7T port map(CN => lbl0_n_541, CP => CTS_20, D => lbl0_n_35, Q => lbl0_counter_busy_counter_state(0));
  lbl0_counter_unsigned_busy_count_reg_1 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN279_lbl0_n_37, Q => lbl0_busy_count(1));
  lbl0_counter_unsigned_busy_count_reg_5 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN274_lbl0_n_38, Q => lbl0_busy_count(5));
  lbl0_counter_unsigned_busy_count_reg_0 : DFXQD1BWP7T port map(CP => CTS_20, DA => lbl0_n_27, DB => lbl0_n_14, Q => lbl0_busy_count(0), SA => FE_PHN315_lbl0_busy_count_0);
  lbl0_g8610 : ND3D0BWP7T port map(A1 => FE_PHN309_lbl0_n_539, A2 => lbl0_n_36, A3 => lbl0_n_21, ZN => lbl0_n_47);
  lbl0_g8611 : OAI211D1BWP7T port map(A1 => lbl0_n_9, A2 => lbl0_n_25, B => lbl0_n_22, C => lbl0_n_17, ZN => lbl0_n_46);
  lbl0_g8612 : OAI32D1BWP7T port map(A1 => lbl0_busy_count(2), A2 => lbl0_n_437, A3 => lbl0_n_15, B1 => lbl0_n_4, B2 => lbl0_n_30, ZN => lbl0_n_45);
  lbl0_g8613 : OAI32D1BWP7T port map(A1 => lbl0_busy_count(4), A2 => lbl0_n_436, A3 => lbl0_n_15, B1 => lbl0_n_2, B2 => lbl0_n_32, ZN => lbl0_n_44);
  lbl0_g8614 : AO22D0BWP7T port map(A1 => lbl0_n_33, A2 => lbl0_busy_count(6), B1 => lbl0_n_24, B2 => lbl0_n_14, Z => lbl0_n_43);
  lbl0_g8615 : AO22D0BWP7T port map(A1 => lbl0_n_31, A2 => lbl0_busy_count(3), B1 => lbl0_n_23, B2 => lbl0_n_14, Z => lbl0_n_42);
  lbl0_g8616 : IOA21D1BWP7T port map(A1 => lbl0_n_446, A2 => FE_DBTN24_rst, B => lbl0_n_36, ZN => lbl0_n_41);
  lbl0_g8617 : AOI32D1BWP7T port map(A1 => memory_ready, A2 => lbl0_n_16, A3 => FE_PHN314_lbl0_mem_com_state_0, B1 => lbl0_n_450, B2 => FE_DBTN24_rst, ZN => lbl0_n_40);
  lbl0_g8620 : MOAI22D0BWP7T port map(A1 => lbl0_n_15, A2 => lbl0_n_12, B1 => lbl0_n_27, B2 => lbl0_busy_count(5), ZN => lbl0_n_38);
  lbl0_g8621 : MOAI22D0BWP7T port map(A1 => lbl0_n_15, A2 => lbl0_n_13, B1 => lbl0_n_27, B2 => lbl0_busy_count(1), ZN => lbl0_n_37);
  lbl0_g8622 : ND2D1BWP7T port map(A1 => lbl0_n_27, A2 => busy, ZN => lbl0_n_35);
  lbl0_g8623 : IOA21D1BWP7T port map(A1 => lbl0_n_20, A2 => busy, B => lbl0_n_18, ZN => lbl0_n_34);
  lbl0_g8624 : IND3D1BWP7T port map(A1 => lbl0_mem_com_state(0), B1 => FE_PHN262_lbl0_mem_com_state_3, B2 => lbl0_n_19, ZN => lbl0_n_36);
  lbl0_g8625 : INVD0BWP7T port map(I => lbl0_n_32, ZN => lbl0_n_33);
  lbl0_g8626 : INVD0BWP7T port map(I => lbl0_n_30, ZN => lbl0_n_31);
  lbl0_g8627 : ND3D0BWP7T port map(A1 => lbl0_n_11, A2 => lbl0_state(2), A3 => lbl0_state(3), ZN => lbl0_n_28);
  lbl0_g8628 : AOI21D0BWP7T port map(A1 => lbl0_n_14, A2 => lbl0_n_436, B => lbl0_n_27, ZN => lbl0_n_32);
  lbl0_g8629 : AOI21D0BWP7T port map(A1 => lbl0_n_14, A2 => lbl0_n_437, B => lbl0_n_27, ZN => lbl0_n_30);
  lbl0_g8632 : IND2D1BWP7T port map(A1 => lbl0_n_20, B1 => lbl0_n_18, ZN => lbl0_n_27);
  lbl0_g8633 : AOI31D0BWP7T port map(A1 => lbl0_n_461, A2 => lbl0_n_5, A3 => lbl0_state(3), B => lbl0_n_532, ZN => lbl0_n_25);
  lbl0_g8634 : OAI32D1BWP7T port map(A1 => lbl0_busy_count(6), A2 => lbl0_n_7, A3 => lbl0_n_436, B1 => lbl0_n_1, B2 => lbl0_n_438, ZN => lbl0_n_24);
  lbl0_g8635 : OAI32D1BWP7T port map(A1 => lbl0_busy_count(3), A2 => lbl0_n_4, A3 => lbl0_n_437, B1 => lbl0_busy_count(2), B2 => lbl0_n_0, ZN => lbl0_n_23);
  lbl0_g8637 : ND2D0BWP7T port map(A1 => clear_memory, A2 => lbl0_n_10, ZN => lbl0_n_21);
  lbl0_g8640 : IND2D1BWP7T port map(A1 => lbl0_n_9, B1 => lbl0_n_536, ZN => lbl0_n_22);
  lbl0_g8643 : INVD0BWP7T port map(I => lbl0_n_17, ZN => lbl0_n_16);
  lbl0_g8644 : INVD1BWP7T port map(I => lbl0_n_15, ZN => lbl0_n_14);
  lbl0_g8645 : XNR2D1BWP7T port map(A1 => FE_PHN258_lbl0_busy_count_0, A2 => lbl0_busy_count(1), ZN => lbl0_n_13);
  lbl0_g8646 : MAOI22D0BWP7T port map(A1 => lbl0_n_439, A2 => lbl0_busy_count(5), B1 => lbl0_n_439, B2 => lbl0_busy_count(5), ZN => lbl0_n_12);
  lbl0_g8647 : CKXOR2D0BWP7T port map(A1 => lbl0_state(1), A2 => lbl0_state(0), Z => lbl0_n_11);
  lbl0_g8648 : AN3D0BWP7T port map(A1 => lbl0_n_541, A2 => lbl0_n_6, A3 => FE_PHN182_lbl0_counter_busy_counter_state_0, Z => lbl0_n_20);
  lbl0_g8649 : NR3D0BWP7T port map(A1 => lbl0_mem_com_state(1), A2 => lbl0_mem_com_state(2), A3 => FE_OFN1_rst, ZN => lbl0_n_19);
  lbl0_g8650 : IND3D1BWP7T port map(A1 => FE_PHN182_lbl0_counter_busy_counter_state_0, B1 => lbl0_counter_busy_counter_state(1), B2 => lbl0_n_541, ZN => lbl0_n_18);
  lbl0_g8651 : IND3D1BWP7T port map(A1 => lbl0_mem_com_state(1), B1 => FE_PHN333_lbl0_mem_com_state_2, B2 => lbl0_n_10, ZN => lbl0_n_17);
  lbl0_g8652 : ND3D0BWP7T port map(A1 => lbl0_n_541, A2 => FE_PHN182_lbl0_counter_busy_counter_state_0, A3 => lbl0_counter_busy_counter_state(1), ZN => lbl0_n_15);
  lbl0_g8653 : NR2XD0BWP7T port map(A1 => FE_PHN262_lbl0_mem_com_state_3, A2 => FE_OFN1_rst, ZN => lbl0_n_10);
  lbl0_g8654 : ND2D1BWP7T port map(A1 => lbl0_mem_com_n_166, A2 => FE_DBTN24_rst, ZN => lbl0_n_9);
  lbl0_g8656 : INVD0BWP7T port map(I => lbl0_n_438, ZN => lbl0_n_7);
  lbl0_mem_com_state_reg_1 : DFD1BWP7T port map(CP => CTS_20, D => lbl0_n_48, Q => FE_PHN256_lbl0_mem_com_state_1, QN => lbl0_n_79);
  lbl0_counter_unsigned_busy_count_reg_4 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN268_lbl0_n_44, Q => lbl0_busy_count(4), QN => lbl0_n_2);
  lbl0_mem_com_state_reg_0 : DFD1BWP7T port map(CP => CTS_20, D => lbl0_n_50, Q => FE_PHN266_lbl0_mem_com_state_0, QN => lbl0_n_67);
  lbl0_mem_com_state_reg_2 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN307_lbl0_n_46, Q => lbl0_mem_com_state(2), QN => lbl0_n_66);
  lbl0_state_reg_1 : DFKCND1BWP7T port map(CN => lbl0_new_state(1), CP => CTS_20, D => FE_DBTN24_rst, Q => lbl0_state(1), QN => lbl0_n_60);
  lbl0_state_reg_4 : DFKCND1BWP7T port map(CN => lbl0_new_state(4), CP => CTS_20, D => FE_DBTN24_rst, Q => lbl0_state(4), QN => lbl0_n_59);
  lbl0_state_reg_3 : DFKCND1BWP7T port map(CN => lbl0_new_state(3), CP => CTS_20, D => FE_DBTN24_rst, Q => lbl0_state(3), QN => lbl0_n_58);
  lbl0_state_reg_2 : DFKCND1BWP7T port map(CN => lbl0_new_state(2), CP => CTS_20, D => FE_DBTN24_rst, Q => lbl0_state(2), QN => lbl0_n_5);
  lbl0_state_reg_0 : DFKCND1BWP7T port map(CN => lbl0_new_state(0), CP => CTS_20, D => FE_DBTN24_rst, Q => lbl0_state(0), QN => lbl0_n_56);
  lbl0_counter_busy_counter_state_reg_1 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN294_lbl0_n_34, Q => FE_PHN164_lbl0_counter_busy_counter_state_1, QN => lbl0_n_6);
  lbl0_counter_unsigned_busy_count_reg_6 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN276_lbl0_n_43, Q => lbl0_busy_count(6), QN => lbl0_n_1);
  lbl0_counter_unsigned_busy_count_reg_3 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN272_lbl0_n_42, Q => lbl0_busy_count(3), QN => lbl0_n_0);
  lbl0_counter_unsigned_busy_count_reg_2 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN269_lbl0_n_45, Q => lbl0_busy_count(2), QN => lbl0_n_4);
  lbl0_g18955 : IND3D1BWP7T port map(A1 => lbl0_n_128, B1 => lbl0_n_536, B2 => lbl0_n_19, ZN => lbl0_n_539);
  lbl0_g18956 : AO222D0BWP7T port map(A1 => lbl0_n_288, A2 => lbl0_n_150, B1 => lbl0_n_317, B2 => lbl0_read_data_reg(6), C1 => lbl0_n_292, C2 => lbl0_n_147, Z => write_memory(6));
  lbl0_g18957 : IAO21D0BWP7T port map(A1 => lbl0_n_164, A2 => lbl0_state(0), B => FE_OFN1_rst, ZN => lbl0_n_541);
  lbl0_g18958 : MAOI22D0BWP7T port map(A1 => lbl0_mem_com_n_175, A2 => lbl0_n_10, B1 => memory_ready, B2 => lbl0_n_17, ZN => lbl0_n_542);
  lbl0_reg_pos0_q_reg_2 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_position_0(2), E => lbl0_e_position_0, Q => position_0(2));
  lbl0_reg_pos0_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_21, D => lbl0_d_position_0(1), E => lbl0_e_position_0, Q => position_0(1));
  lbl0_reg_pos0_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_440, E => lbl0_e_position_0, Q => position_0(0));
  lbl0_reg_pos0_q_reg_7 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_position_0(7), E => lbl0_e_position_0, Q => position_0(7));
  lbl0_reg_pos0_q_reg_8 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_position_0(8), E => lbl0_e_position_0, Q => position_0(8));
  lbl0_reg_pos0_q_reg_4 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_441, E => lbl0_e_position_0, Q => position_0(4));
  lbl0_reg_pos0_q_reg_3 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_position_0(3), E => lbl0_e_position_0, Q => position_0(3));
  lbl0_reg_pos0_q_reg_9 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_443, E => lbl0_e_position_0, Q => position_0(9));
  lbl0_reg_pos0_q_reg_5 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_442, E => lbl0_e_position_0, Q => position_0(5));
  lbl0_reg_pos0_q_reg_6 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_position_0(6), E => lbl0_e_position_0, Q => position_0(6));
  lbl0_reg_n_layer_1_q_reg : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_499, E => lbl0_n_530, Q => lbl0_next_layer_1);
  lbl0_reg_booster_sync_q_reg : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_booster_sync, E => lbl0_n_456, Q => lbl0_booster_sync);
  lbl0_reg_pos1_q_reg_2 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_position_1(2), E => lbl0_e_position_1, Q => position_1(2));
  lbl0_reg_pos1_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_position_1(1), E => lbl0_e_position_1, Q => position_1(1));
  lbl0_reg_pos1_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_position_1(0), E => lbl0_e_position_1, Q => position_1(0));
  lbl0_reg_pos1_q_reg_7 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_21, D => lbl0_d_position_1(7), E => lbl0_e_position_1, Q => position_1(7));
  lbl0_reg_pos1_q_reg_8 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_21, D => lbl0_d_position_1(8), E => lbl0_e_position_1, Q => position_1(8));
  lbl0_reg_pos1_q_reg_4 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_position_1(4), E => lbl0_e_position_1, Q => position_1(4));
  lbl0_reg_pos1_q_reg_3 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_position_1(3), E => lbl0_e_position_1, Q => position_1(3));
  lbl0_reg_pos1_q_reg_9 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_position_1(9), E => lbl0_e_position_1, Q => position_1(9));
  lbl0_reg_pos1_q_reg_5 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_position_1(5), E => lbl0_e_position_1, Q => position_1(5));
  lbl0_reg_pos1_q_reg_6 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_21, D => lbl0_d_position_1(6), E => lbl0_e_position_1, Q => position_1(6));
  lbl0_reg_border_0_q_reg : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_498, E => lbl0_n_531, Q => lbl0_border_0);
  lbl0_reg_border_1_q_reg : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_497, E => lbl0_n_530, Q => lbl0_border_1);
  lbl0_reg_dir_0_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_direction_0(0), E => lbl0_n_457, Q => direction_0(0));
  lbl0_reg_dir_0_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_direction_0(1), E => lbl0_n_457, Q => direction_0(1));
  lbl0_reg_p_state_0_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_448, E => lbl0_n_445, Q => player_state_0(0));
  lbl0_reg_p_state_0_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_449, E => lbl0_n_445, Q => player_state_0(1));
  lbl0_reg_dir_1_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_direction_1(0), E => lbl0_n_457, Q => direction_1(0));
  lbl0_reg_dir_1_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_direction_1(1), E => lbl0_n_457, Q => direction_1(1));
  lbl0_reg_speed_select_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN24_rst, CP => CTS_20, D => lbl0_d_speed_select(0), E => lbl0_n_535, Q => lbl0_n_503);
  lbl0_reg_speed_select_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN24_rst, CP => CTS_20, D => lbl0_d_speed_select(1), E => lbl0_n_535, Q => lbl0_n_502);
  lbl0_reg_p_state_1_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_447, E => lbl0_n_444, Q => player_state_1(0));
  lbl0_reg_p_state_1_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_449, E => lbl0_n_444, Q => player_state_1(1));
  lbl0_reg_boost_audio_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_453, E => lbl0_n_533, Q => boost_audio_0);
  lbl0_reg_boost_audio_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_454, E => lbl0_n_533, Q => boost_audio_1);
  lbl0_reg_n_dir_0_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_next_direction_0(0), E => lbl0_n_452, Q => lbl0_next_direction_0(0));
  lbl0_reg_n_dir_0_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_next_direction_0(1), E => lbl0_n_452, Q => lbl0_next_direction_0(1));
  lbl0_reg_n_dir_1_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_next_direction_1(0), E => lbl0_n_451, Q => lbl0_next_direction_1(0));
  lbl0_reg_n_dir_1_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_next_direction_1(1), E => lbl0_n_451, Q => lbl0_next_direction_1(1));
  lbl0_reg_layer_0_q_reg : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_layer_0, E => lbl0_e_position_0, Q => position_0(10));
  lbl0_reg_layer_1_q_reg : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_layer_1, E => lbl0_e_position_1, Q => position_1(10));
  lbl0_reg_map_select_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_map_select(0), E => lbl0_n_535, Q => map_selected(0));
  lbl0_reg_map_select_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_map_select(1), E => lbl0_n_535, Q => map_selected(1));
  lbl0_reg_move_0_q_reg : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_move_0, E => lbl0_n_456, Q => lbl0_move_0);
  lbl0_reg_r_mem_0_q_reg_3 : EDFKCNQD1BWP7T port map(CN => FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_read_data_reg(3), E => lbl0_n_455, Q => lbl0_read_data_reg(3));
  lbl0_reg_r_mem_0_q_reg_2 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_read_data_reg(2), E => lbl0_n_455, Q => lbl0_read_data_reg(2));
  lbl0_reg_r_mem_0_q_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_read_data_reg(0), E => lbl0_n_455, Q => lbl0_read_data_reg(0));
  lbl0_reg_r_mem_0_q_reg_4 : EDFKCNQD1BWP7T port map(CN => FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_read_data_reg(4), E => lbl0_n_455, Q => lbl0_read_data_reg(4));
  lbl0_reg_r_mem_0_q_reg_6 : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_read_data_reg(6), E => lbl0_n_455, Q => lbl0_read_data_reg(6));
  lbl0_reg_r_mem_0_q_reg_5 : EDFKCNQD1BWP7T port map(CN => FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_read_data_reg(5), E => lbl0_n_455, Q => lbl0_read_data_reg(5));
  lbl0_reg_r_mem_0_q_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_read_data_reg(1), E => lbl0_n_455, Q => lbl0_read_data_reg(1));
  lbl0_reg_r_mem_0_q_reg_7 : EDFKCNQD1BWP7T port map(CN => FE_DBTN24_rst, CP => CTS_20, D => lbl0_d_read_data_reg(7), E => lbl0_n_455, Q => lbl0_read_data_reg(7));
  lbl0_reg_move_1_q_reg : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_d_move_1, E => lbl0_n_456, Q => lbl0_move_1);
  lbl1_g22 : OR3D4BWP7T port map(A1 => lbl1_x_incr3, A2 => lbl1_x_incr2, A3 => lbl1_x_incr1, Z => x_increment_out);
  lbl1_g21 : OR3D4BWP7T port map(A1 => lbl1_y_incr3, A2 => lbl1_y_incr2, A3 => lbl1_y_incr1, Z => y_increment_out);
  lbl1_g18 : CKAN2D8BWP7T port map(A1 => lbl1_we_clr, A2 => lbl1_we_rw, Z => write_enable_out);
  lbl1_g12 : OR2D1BWP7T port map(A1 => lbl1_me_rw, A2 => lbl1_me_clr, Z => FE_OFN4_memory_enable_out);
  lbl1_g23 : CKAN2D1BWP7T port map(A1 => lbl1_ready_rw, A2 => lbl1_ready_clr, Z => memory_ready);
  lbl1_g26 : OR4D4BWP7T port map(A1 => FE_OFN1_rst, A2 => lbl1_clr_rst, A3 => lbl1_rw_rst, A4 => reset_vga_mem, Z => memory_reset_out);
  lbl1_cy_count_reg_4 : DFKCNQD1BWP7T port map(CN => FE_PHN310_lbl1_cy_n_10, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => y_address(4));
  lbl1_cy_count_reg_3 : DFKCNQD1BWP7T port map(CN => lbl1_cy_n_9, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => y_address(3));
  lbl1_cy_g92 : MOAI22D0BWP7T port map(A1 => lbl1_cy_n_8, A2 => y_address(4), B1 => lbl1_cy_n_8, B2 => y_address(4), ZN => lbl1_cy_n_10);
  lbl1_cy_count_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN302_lbl1_cy_n_7, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => y_address(2));
  lbl1_cy_g94 : MOAI22D0BWP7T port map(A1 => lbl1_cy_n_6, A2 => FE_PHN247_y_address_3, B1 => lbl1_cy_n_6, B2 => FE_PHN247_y_address_3, ZN => lbl1_cy_n_9);
  lbl1_cy_g95 : IND2D1BWP7T port map(A1 => lbl1_cy_n_6, B1 => FE_PHN247_y_address_3, ZN => lbl1_cy_n_8);
  lbl1_cy_count_reg_1 : DFKCNQD1BWP7T port map(CN => FE_PHN301_lbl1_cy_n_5, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => y_address(1));
  lbl1_cy_g97 : MOAI22D0BWP7T port map(A1 => lbl1_cy_n_4, A2 => y_address(2), B1 => lbl1_cy_n_4, B2 => y_address(2), ZN => lbl1_cy_n_7);
  lbl1_cy_g98 : IND2D1BWP7T port map(A1 => lbl1_cy_n_4, B1 => y_address(2), ZN => lbl1_cy_n_6);
  lbl1_cy_count_reg_0 : DFKCNQD1BWP7T port map(CN => FE_PHN305_lbl1_cy_n_3, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => y_address(0));
  lbl1_cy_g100 : MOAI22D0BWP7T port map(A1 => lbl1_cy_n_2, A2 => y_address(1), B1 => lbl1_cy_n_2, B2 => y_address(1), ZN => lbl1_cy_n_5);
  lbl1_cy_g101 : IND2D1BWP7T port map(A1 => lbl1_cy_n_2, B1 => y_address(1), ZN => lbl1_cy_n_4);
  lbl1_cy_g102 : MOAI22D0BWP7T port map(A1 => lbl1_cy_n_1, A2 => FE_PHN324_y_address_0, B1 => lbl1_cy_n_1, B2 => y_address(0), ZN => lbl1_cy_n_3);
  lbl1_cy_g103 : IND2D1BWP7T port map(A1 => lbl1_cy_n_1, B1 => y_address(0), ZN => lbl1_cy_n_2);
  lbl1_cy_g104 : ND2D1BWP7T port map(A1 => y_increment_out, A2 => lbl1_cy_prev_incr, ZN => lbl1_cy_n_1);
  lbl1_cy_prev_incr_reg : DFD1BWP7T port map(CP => CTS_18, D => y_increment_out, Q => UNCONNECTED7, QN => lbl1_cy_prev_incr);
  lbl1_cm_g500 : AO221D0BWP7T port map(A1 => lbl1_cm_n_38, A2 => lbl1_cm_n_27, B1 => lbl1_cm_n_28, B2 => lbl1_cm_state(3), C => lbl1_x_incr3, Z => lbl1_we_clr);
  lbl1_cm_g501 : AO31D1BWP7T port map(A1 => lbl1_cm_n_27, A2 => lbl1_cm_n_30, A3 => lbl1_cm_state(0), B => lbl1_cm_state(4), Z => lbl1_clr_rst);
  lbl1_cm_g502 : INR4D0BWP7T port map(A1 => lbl1_cm_n_27, B1 => lbl1_cm_state(1), B2 => lbl1_cm_state(0), B3 => lbl1_cm_state(4), ZN => lbl1_ready_clr);
  lbl1_cm_g503 : CKAN2D1BWP7T port map(A1 => lbl1_x_incr3, A2 => lbl1_cm_state(1), Z => lbl1_y_incr3);
  lbl1_cm_g504 : CKND1BWP7T port map(I => lbl1_cm_n_38, ZN => lbl1_cm_n_28);
  lbl1_cm_g505 : NR2XD0BWP7T port map(A1 => lbl1_cm_n_30, A2 => lbl1_cm_state(2), ZN => lbl1_me_clr);
  lbl1_cm_g506 : ND2D1BWP7T port map(A1 => lbl1_cm_state(0), A2 => lbl1_cm_state(1), ZN => lbl1_cm_n_38);
  lbl1_cm_g507 : INR2D1BWP7T port map(A1 => lbl1_cm_state(0), B1 => lbl1_cm_state(3), ZN => lbl1_cm_n_364_BAR);
  lbl1_cm_g508 : NR2XD0BWP7T port map(A1 => lbl1_cm_n_29, A2 => lbl1_cm_n_31, ZN => lbl1_x_incr3);
  lbl1_cm_g509 : NR2XD0BWP7T port map(A1 => lbl1_cm_state(2), A2 => lbl1_cm_state(3), ZN => lbl1_cm_n_27);
  lbl1_cm_g852 : OAI21D0BWP7T port map(A1 => lbl1_cm_n_3, A2 => lbl1_cm_n_22, B => lbl1_cm_n_21, ZN => lbl1_cm_n_26);
  lbl1_cm_g853 : IOA21D1BWP7T port map(A1 => lbl1_cm_n_2, A2 => lbl1_cm_n_52, B => lbl1_cm_n_21, ZN => lbl1_cm_n_25);
  lbl1_cm_state_reg_4 : DFKCNQD1BWP7T port map(CN => lbl1_cm_n_14, CP => CTS_18, D => lbl1_cm_n_19, Q => lbl1_cm_state(4));
  lbl1_cm_g855 : OAI22D0BWP7T port map(A1 => lbl1_cm_n_54, A2 => FE_PHN339_lbl1_cm_state_0, B1 => lbl1_cm_n_5, B2 => FE_OFN1_rst, ZN => lbl1_cm_n_24);
  lbl1_cm_g856 : AO32D1BWP7T port map(A1 => lbl1_cm_n_2, A2 => lbl1_cm_n_12, A3 => lbl1_cm_n_8, B1 => lbl1_cm_n_19, B2 => lbl1_cm_n_13, Z => lbl1_cm_n_23);
  lbl1_cm_g857 : AOI211XD0BWP7T port map(A1 => lbl1_cm_n_4, A2 => lbl1_cm_n_38, B => lbl1_cm_n_53, C => lbl1_cm_n_55, ZN => FE_PHN156_lbl1_cm_n_22);
  lbl1_cm_g859 : OAI21D0BWP7T port map(A1 => lbl1_cm_n_15, A2 => lbl1_cm_n_13, B => lbl1_cm_n_16, ZN => lbl1_cm_n_21);
  lbl1_cm_g860 : INR2D1BWP7T port map(A1 => lbl1_cm_n_16, B1 => lbl1_cm_n_15, ZN => lbl1_cm_n_19);
  lbl1_cm_g863 : NR2XD0BWP7T port map(A1 => lbl1_cm_n_12, A2 => FE_OFN1_rst, ZN => lbl1_cm_n_16);
  lbl1_cm_g864 : INVD0BWP7T port map(I => lbl1_cm_n_13, ZN => lbl1_cm_n_14);
  lbl1_cm_g865 : IND4D0BWP7T port map(A1 => lbl1_cm_n_1, B1 => x_address(3), B2 => x_address(0), B3 => x_address(2), ZN => lbl1_cm_n_15);
  lbl1_cm_g866 : IND4D0BWP7T port map(A1 => lbl1_cm_n_6, B1 => y_address(2), B2 => y_address(1), B3 => y_address(4), ZN => lbl1_cm_n_13);
  lbl1_cm_g867 : ND2D0BWP7T port map(A1 => lbl1_cm_n_7, A2 => lbl1_cm_n_31, ZN => lbl1_cm_n_11);
  lbl1_cm_g868 : IND2D1BWP7T port map(A1 => lbl1_cm_n_31, B1 => lbl1_cm_n_7, ZN => lbl1_cm_n_12);
  lbl1_cm_g870 : OA21D0BWP7T port map(A1 => lbl1_cm_state(1), A2 => lbl1_cm_state(3), B => lbl1_cm_state(0), Z => lbl1_cm_n_9);
  lbl1_cm_g871 : OAI22D0BWP7T port map(A1 => lbl1_cm_n_364_BAR, A2 => lbl1_cm_n_30, B1 => lbl1_cm_n_0, B2 => lbl1_cm_state(1), ZN => FE_PHN343_lbl1_cm_n_8);
  lbl1_cm_g872 : ND2D0BWP7T port map(A1 => y_address(0), A2 => FE_PHN247_y_address_3, ZN => lbl1_cm_n_6);
  lbl1_cm_g873 : ND2D1BWP7T port map(A1 => lbl1_ready_clr, A2 => clear_memory, ZN => lbl1_cm_n_5);
  lbl1_cm_g874 : NR2XD0BWP7T port map(A1 => lbl1_cm_n_38, A2 => lbl1_cm_state(2), ZN => lbl1_cm_n_7);
  lbl1_cm_g875 : INVD0BWP7T port map(I => lbl1_cm_n_2, ZN => lbl1_cm_n_3);
  lbl1_cm_g876 : ND2D0BWP7T port map(A1 => x_address(1), A2 => x_address(4), ZN => lbl1_cm_n_1);
  lbl1_cm_g877 : NR2D1BWP7T port map(A1 => lbl1_cm_n_31, A2 => lbl1_cm_state(2), ZN => lbl1_cm_n_4);
  lbl1_cm_g878 : NR2XD0BWP7T port map(A1 => lbl1_ready_clr, A2 => FE_OFN1_rst, ZN => lbl1_cm_n_2);
  lbl1_cm_g2 : OAI21D0BWP7T port map(A1 => lbl1_cm_n_29, A2 => lbl1_cm_n_9, B => lbl1_cm_n_11, ZN => FE_PHN174_lbl1_cm_n_52);
  lbl1_cm_g887 : NR3D0BWP7T port map(A1 => lbl1_cm_n_38, A2 => lbl1_cm_n_29, A3 => lbl1_cm_state(3), ZN => lbl1_cm_n_53);
  lbl1_cm_g888 : IND2D1BWP7T port map(A1 => lbl1_cm_state(4), B1 => lbl1_cm_n_2, ZN => lbl1_cm_n_54);
  lbl1_cm_g889 : NR2D1BWP7T port map(A1 => lbl1_cm_state(0), A2 => lbl1_cm_n_31, ZN => lbl1_cm_n_55);
  lbl1_cm_state_reg_3 : DFD1BWP7T port map(CP => CTS_20, D => lbl1_cm_n_26, Q => lbl1_cm_state(3), QN => lbl1_cm_n_31);
  lbl1_cm_state_reg_2 : DFD1BWP7T port map(CP => CTS_20, D => lbl1_cm_n_25, Q => lbl1_cm_state(2), QN => lbl1_cm_n_29);
  lbl1_cm_state_reg_1 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN308_lbl1_cm_n_23, Q => lbl1_cm_state(1), QN => lbl1_cm_n_30);
  lbl1_cm_state_reg_0 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN293_lbl1_cm_n_24, Q => lbl1_cm_state(0), QN => lbl1_cm_n_0);
  lbl1_cex_g175 : OR2D1BWP7T port map(A1 => lbl1_cex_n_5, A2 => lbl1_cex_n_4, Z => lbl1_x_incr2);
  lbl1_cex_g176 : INR2XD0BWP7T port map(A1 => lbl1_cex_state(1), B1 => lbl1_cex_state(0), ZN => lbl1_cex_n_4);
  lbl1_cex_g177 : INR2XD0BWP7T port map(A1 => lbl1_cex_state(0), B1 => lbl1_cex_state(1), ZN => lbl1_cex_n_5);
  lbl1_cex_state_reg_0 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN304_lbl1_cex_n_3, Q => lbl1_cex_state(0));
  lbl1_cex_state_reg_1 : DFQD1BWP7T port map(CP => CTS_20, D => lbl1_cex_n_2, Q => lbl1_cex_state(1));
  lbl1_cex_g145 : IAO21D0BWP7T port map(A1 => lbl1_cex_n_0, A2 => FE_PHN157_lbl1_cex_n_4, B => FE_OFN1_rst, ZN => lbl1_cex_n_3);
  lbl1_cex_g146 : NR2XD0BWP7T port map(A1 => FE_PHN275_lbl1_cex_n_1, A2 => FE_OFN1_rst, ZN => lbl1_cex_n_2);
  lbl1_cex_g147 : AOI21D0BWP7T port map(A1 => x_increment, A2 => lbl1_cex_state(0), B => lbl1_x_incr2, ZN => lbl1_cex_n_1);
  lbl1_cex_g148 : INR2D1BWP7T port map(A1 => x_increment, B1 => lbl1_cex_n_5, ZN => lbl1_cex_n_0);
  lbl1_rw_g1132 : AN2D1BWP7T port map(A1 => lbl1_rw_n_79, A2 => lbl1_rw_n_87, Z => lbl1_ready_rw);
  lbl1_rw_g1133 : CKAN2D1BWP7T port map(A1 => lbl1_rw_n_79, A2 => lbl1_rw_state(0), Z => lbl1_rw_rst);
  lbl1_rw_g1134 : OAI21D0BWP7T port map(A1 => lbl1_rw_n_78, A2 => lbl1_rw_n_97, B => lbl1_rw_n_84, ZN => lbl1_me_rw);
  lbl1_rw_g1135 : OAI221D0BWP7T port map(A1 => lbl1_rw_n_74, A2 => lbl1_rw_n_80, B1 => lbl1_rw_n_85, B2 => lbl1_rw_n_81, C => lbl1_rw_n_76, ZN => lbl1_y_incr1);
  lbl1_rw_g1136 : NR4D0BWP7T port map(A1 => lbl1_rw_n_74, A2 => lbl1_rw_state(3), A3 => lbl1_rw_state(4), A4 => lbl1_rw_state(5), ZN => lbl1_rw_n_79);
  lbl1_rw_g1137 : OAI221D0BWP7T port map(A1 => lbl1_rw_n_96, A2 => lbl1_rw_state(4), B1 => lbl1_rw_state(1), B2 => lbl1_rw_n_80, C => lbl1_rw_n_76, ZN => lbl1_x_incr1);
  lbl1_rw_g1138 : MOAI22D0BWP7T port map(A1 => lbl1_rw_n_75, A2 => lbl1_rw_n_87, B1 => lbl1_rw_n_97, B2 => lbl1_rw_n_84, ZN => lbl1_we_rw);
  lbl1_rw_g1139 : ND2D5BWP7T port map(A1 => lbl1_rw_n_76, A2 => lbl1_rw_n_77, ZN => w_increment_out);
  lbl1_rw_g1140 : IAO21D0BWP7T port map(A1 => lbl1_rw_n_96, A2 => lbl1_rw_n_87, B => lbl1_rw_n_94, ZN => lbl1_rw_n_78);
  lbl1_rw_g1141 : IND2D1BWP7T port map(A1 => lbl1_rw_n_80, B1 => lbl1_rw_n_74, ZN => lbl1_rw_n_77);
  lbl1_rw_g1142 : NR2XD0BWP7T port map(A1 => lbl1_rw_n_83, A2 => lbl1_rw_n_85, ZN => lbl1_rw_n_94);
  lbl1_rw_g1143 : AN2D0BWP7T port map(A1 => lbl1_rw_n_96, A2 => lbl1_rw_n_84, Z => lbl1_rw_n_75);
  lbl1_rw_g1144 : OR2D1BWP7T port map(A1 => lbl1_rw_n_82, A2 => lbl1_rw_n_74, Z => lbl1_rw_n_76);
  lbl1_rw_g1145 : IND2D1BWP7T port map(A1 => lbl1_rw_state(2), B1 => lbl1_rw_n_85, ZN => lbl1_rw_n_74);
  lbl1_rw_g1146 : IND2D1BWP7T port map(A1 => lbl1_rw_state(4), B1 => lbl1_rw_state(3), ZN => lbl1_rw_n_80);
  lbl1_rw_g1147 : ND2D1BWP7T port map(A1 => lbl1_rw_n_85, A2 => lbl1_rw_state(2), ZN => lbl1_rw_n_96);
  lbl1_rw_g1148 : ND2D1BWP7T port map(A1 => lbl1_rw_n_87, A2 => lbl1_rw_state(2), ZN => lbl1_rw_n_83);
  lbl1_rw_g1149 : IND2D1BWP7T port map(A1 => lbl1_rw_state(4), B1 => lbl1_rw_state(2), ZN => lbl1_rw_n_81);
  lbl1_rw_g1150 : ND2D1BWP7T port map(A1 => lbl1_rw_n_86, A2 => lbl1_rw_state(4), ZN => lbl1_rw_n_82);
  lbl1_rw_g1151 : CKND2D1BWP7T port map(A1 => lbl1_rw_state(4), A2 => lbl1_rw_state(3), ZN => lbl1_rw_n_97);
  lbl1_rw_state_reg_2 : DFQD1BWP7T port map(CP => CTS_20, D => lbl1_rw_n_72, Q => lbl1_rw_state(2));
  lbl1_rw_state_reg_4 : DFQD1BWP7T port map(CP => CTS_20, D => lbl1_rw_n_70, Q => lbl1_rw_state(4));
  lbl1_rw_g2244 : ND2D1BWP7T port map(A1 => lbl1_rw_n_69, A2 => lbl1_rw_n_56, ZN => lbl1_rw_n_73);
  lbl1_rw_g2245 : OR4D1BWP7T port map(A1 => lbl1_rw_n_60, A2 => lbl1_rw_n_62, A3 => lbl1_rw_n_66, A4 => lbl1_rw_n_61, Z => lbl1_rw_n_72);
  lbl1_rw_g2246 : ND3D0BWP7T port map(A1 => lbl1_rw_n_64, A2 => lbl1_rw_n_57, A3 => lbl1_rw_n_50, ZN => lbl1_rw_n_71);
  lbl1_rw_g2248 : OR3D1BWP7T port map(A1 => FE_PHN186_lbl1_rw_n_0, A2 => lbl1_rw_n_65, A3 => lbl1_rw_n_67, Z => lbl1_rw_n_70);
  lbl1_rw_g2249 : AOI211XD0BWP7T port map(A1 => lbl1_rw_n_62, A2 => lbl1_rw_n_38, B => lbl1_rw_n_63, C => lbl1_rw_n_59, ZN => lbl1_rw_n_69);
  lbl1_rw_g2250 : IND3D1BWP7T port map(A1 => lbl1_rw_n_67, B1 => lbl1_rw_n_26, B2 => lbl1_rw_n_53, ZN => lbl1_rw_n_68);
  lbl1_rw_g2251 : OAI221D0BWP7T port map(A1 => lbl1_rw_n_37, A2 => lbl1_rw_n_50, B1 => lbl1_rw_n_47, B2 => lbl1_rw_n_36, C => lbl1_rw_n_43, ZN => lbl1_rw_n_66);
  lbl1_rw_g2252 : OAI22D0BWP7T port map(A1 => lbl1_rw_n_56, A2 => lbl1_rw_n_38, B1 => lbl1_rw_n_36, B2 => lbl1_rw_n_50, ZN => lbl1_rw_n_67);
  lbl1_rw_g2254 : OAI211D1BWP7T port map(A1 => lbl1_rw_n_39, A2 => lbl1_rw_n_55, B => lbl1_rw_n_54, C => lbl1_rw_n_44, ZN => lbl1_rw_n_65);
  lbl1_rw_g2255 : MAOI22D0BWP7T port map(A1 => lbl1_rw_n_41, A2 => FE_PHN152_lbl1_rw_n_27, B1 => lbl1_rw_n_56, B2 => lbl1_rw_n_39, ZN => lbl1_rw_n_64);
  lbl1_rw_g2256 : OAI22D0BWP7T port map(A1 => lbl1_rw_n_55, A2 => lbl1_rw_n_38, B1 => lbl1_rw_n_45, B2 => lbl1_rw_n_3, ZN => lbl1_rw_n_63);
  lbl1_rw_g2257 : NR2D1BWP7T port map(A1 => lbl1_rw_n_56, A2 => lbl1_rw_n_38, ZN => lbl1_rw_n_61);
  lbl1_rw_g2258 : IOA21D1BWP7T port map(A1 => lbl1_rw_n_37, A2 => lbl1_rw_n_51, B => lbl1_rw_n_57, ZN => lbl1_rw_n_62);
  lbl1_rw_g2259 : OAI22D0BWP7T port map(A1 => lbl1_rw_n_46, A2 => lbl1_rw_n_85, B1 => lbl1_rw_n_49, B2 => lbl1_rw_n_81, ZN => lbl1_rw_n_60);
  lbl1_rw_g2260 : OAI22D0BWP7T port map(A1 => lbl1_rw_n_37, A2 => lbl1_rw_n_47, B1 => lbl1_rw_n_49, B2 => lbl1_rw_n_80, ZN => lbl1_rw_n_59);
  lbl1_rw_g2261 : OAI22D0BWP7T port map(A1 => lbl1_rw_n_45, A2 => lbl1_rw_n_4, B1 => lbl1_rw_n_49, B2 => FE_PHN342_lbl1_rw_n_84, ZN => lbl1_rw_n_58);
  lbl1_rw_g2262 : ND2D1BWP7T port map(A1 => lbl1_rw_n_36, A2 => lbl1_rw_n_52, ZN => lbl1_rw_n_57);
  lbl1_rw_g2263 : ND2D1BWP7T port map(A1 => lbl1_rw_n_37, A2 => lbl1_rw_n_52, ZN => lbl1_rw_n_56);
  lbl1_rw_g2264 : AO21D0BWP7T port map(A1 => lbl1_rw_n_85, A2 => lbl1_rw_state(2), B => lbl1_rw_n_45, Z => lbl1_rw_n_54);
  lbl1_rw_g2265 : OAI21D0BWP7T port map(A1 => lbl1_rw_n_96, A2 => lbl1_rw_n_97, B => lbl1_rw_n_48, ZN => lbl1_rw_n_53);
  lbl1_rw_g2266 : ND2D1BWP7T port map(A1 => lbl1_rw_n_36, A2 => lbl1_rw_n_51, ZN => lbl1_rw_n_55);
  lbl1_rw_g2267 : INVD0BWP7T port map(I => lbl1_rw_n_49, ZN => lbl1_rw_n_48);
  lbl1_rw_g2268 : NR2XD0BWP7T port map(A1 => lbl1_rw_n_34, A2 => lbl1_rw_n_42, ZN => lbl1_rw_n_52);
  lbl1_rw_g2269 : NR2D1BWP7T port map(A1 => lbl1_rw_n_35, A2 => lbl1_rw_n_42, ZN => lbl1_rw_n_51);
  lbl1_rw_g2270 : ND2D1BWP7T port map(A1 => lbl1_rw_n_35, A2 => lbl1_rw_n_40, ZN => lbl1_rw_n_50);
  lbl1_rw_g2271 : IND2D1BWP7T port map(A1 => lbl1_rw_state(0), B1 => lbl1_rw_n_41, ZN => lbl1_rw_n_49);
  lbl1_rw_g2272 : CKND1BWP7T port map(I => lbl1_rw_n_0, ZN => lbl1_rw_n_46);
  lbl1_rw_g2273 : OAI21D0BWP7T port map(A1 => lbl1_rw_n_24, A2 => lbl1_rw_n_25, B => lbl1_rw_n_41, ZN => lbl1_rw_n_44);
  lbl1_rw_g2274 : OAI21D0BWP7T port map(A1 => lbl1_rw_n_28, A2 => lbl1_rw_n_94, B => lbl1_rw_n_41, ZN => lbl1_rw_n_43);
  lbl1_rw_g2275 : ND2D1BWP7T port map(A1 => lbl1_rw_n_34, A2 => lbl1_rw_n_40, ZN => lbl1_rw_n_47);
  lbl1_rw_g2277 : IND2D1BWP7T port map(A1 => lbl1_rw_n_97, B1 => lbl1_rw_n_41, ZN => lbl1_rw_n_45);
  lbl1_rw_g2279 : IND3D1BWP7T port map(A1 => FE_OFN1_rst, B1 => lbl1_rw_n_33, B2 => write_enable, ZN => lbl1_rw_n_42);
  lbl1_rw_g2280 : NR3D0BWP7T port map(A1 => lbl1_ready_rw, A2 => lbl1_rw_n_33, A3 => FE_OFN1_rst, ZN => lbl1_rw_n_41);
  lbl1_rw_g2281 : INVD1BWP7T port map(I => lbl1_rw_n_39, ZN => lbl1_rw_n_38);
  lbl1_rw_g2282 : INR3D0BWP7T port map(A1 => lbl1_rw_n_33, B1 => FE_OFN1_rst, B2 => write_enable, ZN => lbl1_rw_n_40);
  lbl1_rw_g2283 : NR4D0BWP7T port map(A1 => lbl1_rw_n_32, A2 => lbl1_rw_n_8, A3 => lbl1_rw_n_29, A4 => lbl1_rw_n_7, ZN => lbl1_rw_n_39);
  lbl1_rw_g2284 : INVD1BWP7T port map(I => lbl1_rw_n_37, ZN => lbl1_rw_n_36);
  lbl1_rw_g2285 : NR4D1BWP7T port map(A1 => lbl1_rw_n_31, A2 => lbl1_rw_n_11, A3 => lbl1_rw_n_15, A4 => lbl1_rw_n_14, ZN => lbl1_rw_n_37);
  lbl1_rw_g2286 : INVD1BWP7T port map(I => lbl1_rw_n_35, ZN => lbl1_rw_n_34);
  lbl1_rw_g2287 : NR4D0BWP7T port map(A1 => lbl1_rw_n_30, A2 => lbl1_rw_n_10, A3 => lbl1_rw_n_9, A4 => lbl1_rw_n_16, ZN => lbl1_rw_n_35);
  lbl1_rw_g2288 : NR4D0BWP7T port map(A1 => lbl1_rw_n_5, A2 => lbl1_rw_n_85, A3 => lbl1_rw_n_87, A4 => lbl1_rw_state(2), ZN => lbl1_rw_n_33);
  lbl1_rw_g2289 : ND4D0BWP7T port map(A1 => lbl1_rw_n_19, A2 => lbl1_rw_n_20, A3 => lbl1_rw_n_22, A4 => lbl1_rw_n_21, ZN => lbl1_rw_n_32);
  lbl1_rw_g2290 : ND2D1BWP7T port map(A1 => lbl1_rw_n_17, A2 => lbl1_rw_n_18, ZN => lbl1_rw_n_31);
  lbl1_rw_g2291 : ND2D1BWP7T port map(A1 => lbl1_rw_n_13, A2 => lbl1_rw_n_12, ZN => lbl1_rw_n_30);
  lbl1_rw_g2292 : ND2D1BWP7T port map(A1 => lbl1_rw_n_6, A2 => lbl1_rw_n_23, ZN => lbl1_rw_n_29);
  lbl1_rw_g2293 : AOI21D0BWP7T port map(A1 => lbl1_rw_n_82, A2 => lbl1_rw_n_1, B => lbl1_rw_n_96, ZN => lbl1_rw_n_28);
  lbl1_rw_g2294 : OAI32D1BWP7T port map(A1 => lbl1_rw_state(1), A2 => lbl1_rw_state(5), A3 => lbl1_rw_n_87, B1 => lbl1_rw_n_85, B2 => lbl1_rw_n_2, ZN => lbl1_rw_n_27);
  lbl1_rw_g2295 : IND3D1BWP7T port map(A1 => FE_OFN1_rst, B1 => go_to, B2 => lbl1_ready_rw, ZN => lbl1_rw_n_26);
  lbl1_rw_g2296 : AOI21D0BWP7T port map(A1 => lbl1_rw_n_83, A2 => lbl1_rw_state(1), B => lbl1_rw_n_82, ZN => lbl1_rw_n_25);
  lbl1_rw_g2297 : AOI21D0BWP7T port map(A1 => lbl1_rw_n_81, A2 => lbl1_rw_n_86, B => lbl1_rw_n_87, ZN => lbl1_rw_n_24);
  lbl1_rw_g2298 : XNR2D1BWP7T port map(A1 => write_memory(6), A2 => lbl1_cur_w(6), ZN => lbl1_rw_n_23);
  lbl1_rw_g2299 : XNR2D1BWP7T port map(A1 => write_memory(3), A2 => lbl1_cur_w(3), ZN => lbl1_rw_n_22);
  lbl1_rw_g2300 : XNR2D1BWP7T port map(A1 => write_memory(2), A2 => FE_PHN212_lbl1_cur_w_2, ZN => lbl1_rw_n_21);
  lbl1_rw_g2301 : XNR2D1BWP7T port map(A1 => write_memory(1), A2 => FE_PHN214_lbl1_cur_w_1, ZN => lbl1_rw_n_20);
  lbl1_rw_g2302 : XNR2D1BWP7T port map(A1 => write_memory(0), A2 => lbl1_cur_w(0), ZN => lbl1_rw_n_19);
  lbl1_rw_g2303 : XNR2D1BWP7T port map(A1 => address(7), A2 => y_address(2), ZN => lbl1_rw_n_18);
  lbl1_rw_g2304 : XNR2D1BWP7T port map(A1 => address(6), A2 => y_address(1), ZN => lbl1_rw_n_17);
  lbl1_rw_g2305 : CKXOR2D1BWP7T port map(A1 => address(0), A2 => x_address(0), Z => lbl1_rw_n_16);
  lbl1_rw_g2306 : CKXOR2D1BWP7T port map(A1 => address(9), A2 => y_address(4), Z => lbl1_rw_n_15);
  lbl1_rw_g2307 : CKXOR2D1BWP7T port map(A1 => address(8), A2 => y_address(3), Z => lbl1_rw_n_14);
  lbl1_rw_g2308 : XNR2D1BWP7T port map(A1 => address(2), A2 => x_address(2), ZN => lbl1_rw_n_13);
  lbl1_rw_g2309 : XNR2D1BWP7T port map(A1 => address(1), A2 => x_address(1), ZN => lbl1_rw_n_12);
  lbl1_rw_g2310 : CKXOR2D1BWP7T port map(A1 => address(5), A2 => y_address(0), Z => lbl1_rw_n_11);
  lbl1_rw_g2311 : CKXOR2D1BWP7T port map(A1 => address(4), A2 => x_address(4), Z => lbl1_rw_n_10);
  lbl1_rw_g2312 : CKXOR2D1BWP7T port map(A1 => address(3), A2 => x_address(3), Z => lbl1_rw_n_9);
  lbl1_rw_g2313 : CKXOR2D1BWP7T port map(A1 => write_memory(5), A2 => lbl1_cur_w(5), Z => lbl1_rw_n_8);
  lbl1_rw_g2314 : CKXOR2D1BWP7T port map(A1 => write_memory(4), A2 => lbl1_cur_w(4), Z => lbl1_rw_n_7);
  lbl1_rw_g2315 : XNR2D1BWP7T port map(A1 => write_memory(7), A2 => lbl1_cur_w(7), ZN => lbl1_rw_n_6);
  lbl1_rw_g2316 : OR2D1BWP7T port map(A1 => lbl1_rw_state(4), A2 => lbl1_rw_state(3), Z => lbl1_rw_n_5);
  lbl1_rw_g2317 : INVD0BWP7T port map(I => lbl1_rw_n_3, ZN => lbl1_rw_n_4);
  lbl1_rw_g2318 : INVD0BWP7T port map(I => lbl1_rw_n_1, ZN => lbl1_rw_n_2);
  lbl1_rw_g2319 : INR2D1BWP7T port map(A1 => lbl1_rw_n_87, B1 => lbl1_rw_n_96, ZN => lbl1_rw_n_3);
  lbl1_rw_g2320 : CKND2D1BWP7T port map(A1 => lbl1_rw_state(0), A2 => lbl1_rw_state(4), ZN => lbl1_rw_n_1);
  lbl1_rw_g2 : INR3D0BWP7T port map(A1 => lbl1_rw_n_41, B1 => lbl1_rw_n_1, B2 => lbl1_rw_state(2), ZN => lbl1_rw_n_0);
  lbl1_rw_state_reg_3 : DFD1BWP7T port map(CP => CTS_20, D => lbl1_rw_n_73, Q => lbl1_rw_state(3), QN => lbl1_rw_n_86);
  lbl1_rw_state_reg_5 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN149_lbl1_rw_n_58, Q => lbl1_rw_state(5), QN => lbl1_rw_n_84);
  lbl1_rw_state_reg_0 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN291_lbl1_rw_n_68, Q => lbl1_rw_state(0), QN => lbl1_rw_n_87);
  lbl1_rw_state_reg_1 : DFD1BWP7T port map(CP => CTS_20, D => lbl1_rw_n_71, Q => lbl1_rw_state(1), QN => lbl1_rw_n_85);
  lbl1_cey_g175 : OR2D1BWP7T port map(A1 => lbl1_cey_n_5, A2 => lbl1_cey_n_4, Z => lbl1_y_incr2);
  lbl1_cey_g176 : INR2XD0BWP7T port map(A1 => lbl1_cey_state(1), B1 => lbl1_cey_state(0), ZN => lbl1_cey_n_4);
  lbl1_cey_g177 : INR2XD0BWP7T port map(A1 => lbl1_cey_state(0), B1 => lbl1_cey_state(1), ZN => lbl1_cey_n_5);
  lbl1_cey_state_reg_0 : DFQD1BWP7T port map(CP => CTS_20, D => lbl1_cey_n_3, Q => lbl1_cey_state(0));
  lbl1_cey_state_reg_1 : DFQD1BWP7T port map(CP => CTS_20, D => lbl1_cey_n_2, Q => lbl1_cey_state(1));
  lbl1_cey_g145 : IAO21D0BWP7T port map(A1 => lbl1_cey_n_0, A2 => FE_PHN154_lbl1_cey_n_4, B => FE_OFN1_rst, ZN => FE_PHN303_lbl1_cey_n_3);
  lbl1_cey_g146 : NR2XD0BWP7T port map(A1 => FE_PHN277_lbl1_cey_n_1, A2 => FE_OFN1_rst, ZN => lbl1_cey_n_2);
  lbl1_cey_g147 : AOI21D0BWP7T port map(A1 => y_increment, A2 => lbl1_cey_state(0), B => lbl1_y_incr2, ZN => lbl1_cey_n_1);
  lbl1_cey_g148 : INR2D1BWP7T port map(A1 => y_increment, B1 => lbl1_cey_n_5, ZN => lbl1_cey_n_0);
  lbl1_cw_count_reg_7 : DFKCNQD1BWP7T port map(CN => FE_PHN297_lbl1_cw_n_16, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => lbl1_cur_w(7));
  lbl1_cw_count_reg_6 : DFKCNQD1BWP7T port map(CN => lbl1_cw_n_15, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => FE_PHN191_lbl1_cur_w_6);
  lbl1_cw_g144 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_14, A2 => lbl1_cur_w(7), B1 => lbl1_cw_n_14, B2 => lbl1_cur_w(7), ZN => lbl1_cw_n_16);
  lbl1_cw_count_reg_5 : DFKCNQD1BWP7T port map(CN => lbl1_cw_n_13, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => FE_PHN326_lbl1_cur_w_5);
  lbl1_cw_g146 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_12, A2 => lbl1_cur_w(6), B1 => lbl1_cw_n_12, B2 => lbl1_cur_w(6), ZN => lbl1_cw_n_15);
  lbl1_cw_g147 : IND2D1BWP7T port map(A1 => lbl1_cw_n_12, B1 => lbl1_cur_w(6), ZN => lbl1_cw_n_14);
  lbl1_cw_count_reg_4 : DFKCNQD1BWP7T port map(CN => lbl1_cw_n_11, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => FE_PHN197_lbl1_cur_w_4);
  lbl1_cw_g149 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_10, A2 => lbl1_cur_w(5), B1 => lbl1_cw_n_10, B2 => lbl1_cur_w(5), ZN => lbl1_cw_n_13);
  lbl1_cw_g150 : IND2D1BWP7T port map(A1 => lbl1_cw_n_10, B1 => lbl1_cur_w(5), ZN => lbl1_cw_n_12);
  lbl1_cw_count_reg_3 : DFKCNQD1BWP7T port map(CN => lbl1_cw_n_9, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => FE_PHN332_lbl1_cur_w_3);
  lbl1_cw_g152 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_8, A2 => lbl1_cur_w(4), B1 => lbl1_cw_n_8, B2 => lbl1_cur_w(4), ZN => lbl1_cw_n_11);
  lbl1_cw_g153 : IND2D1BWP7T port map(A1 => lbl1_cw_n_8, B1 => lbl1_cur_w(4), ZN => lbl1_cw_n_10);
  lbl1_cw_count_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN299_lbl1_cw_n_7, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => lbl1_cur_w(2));
  lbl1_cw_g155 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_6, A2 => lbl1_cur_w(3), B1 => lbl1_cw_n_6, B2 => lbl1_cur_w(3), ZN => lbl1_cw_n_9);
  lbl1_cw_g156 : IND2D1BWP7T port map(A1 => lbl1_cw_n_6, B1 => lbl1_cur_w(3), ZN => lbl1_cw_n_8);
  lbl1_cw_count_reg_1 : DFKCNQD1BWP7T port map(CN => lbl1_cw_n_5, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => lbl1_cur_w(1));
  lbl1_cw_g158 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_4, A2 => FE_PHN212_lbl1_cur_w_2, B1 => lbl1_cw_n_4, B2 => FE_PHN212_lbl1_cur_w_2, ZN => lbl1_cw_n_7);
  lbl1_cw_g159 : IND2D1BWP7T port map(A1 => lbl1_cw_n_4, B1 => FE_PHN212_lbl1_cur_w_2, ZN => lbl1_cw_n_6);
  lbl1_cw_count_reg_0 : DFKCNQD1BWP7T port map(CN => FE_PHN288_lbl1_cw_n_3, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => lbl1_cur_w(0));
  lbl1_cw_g161 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_2, A2 => FE_PHN214_lbl1_cur_w_1, B1 => lbl1_cw_n_2, B2 => FE_PHN214_lbl1_cur_w_1, ZN => lbl1_cw_n_5);
  lbl1_cw_g162 : IND2D1BWP7T port map(A1 => lbl1_cw_n_2, B1 => FE_PHN214_lbl1_cur_w_1, ZN => lbl1_cw_n_4);
  lbl1_cw_g163 : MOAI22D0BWP7T port map(A1 => lbl1_cw_n_1, A2 => FE_PHN200_lbl1_cur_w_0, B1 => lbl1_cw_n_1, B2 => FE_PHN200_lbl1_cur_w_0, ZN => lbl1_cw_n_3);
  lbl1_cw_g164 : IND2D1BWP7T port map(A1 => lbl1_cw_n_1, B1 => FE_PHN200_lbl1_cur_w_0, ZN => lbl1_cw_n_2);
  lbl1_cw_g165 : ND2D1BWP7T port map(A1 => w_increment_out, A2 => lbl1_cw_prev_incr, ZN => lbl1_cw_n_1);
  lbl1_cw_prev_incr_reg : DFD1BWP7T port map(CP => CTS_20, D => w_increment_out, Q => UNCONNECTED8, QN => lbl1_cw_prev_incr);
  lbl1_cx_count_reg_4 : DFKCNQD1BWP7T port map(CN => FE_PHN300_lbl1_cx_n_10, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => x_address(4));
  lbl1_cx_count_reg_3 : DFKCNQD1BWP7T port map(CN => lbl1_cx_n_9, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => FE_PHN257_x_address_3);
  lbl1_cx_g92 : MOAI22D0BWP7T port map(A1 => lbl1_cx_n_8, A2 => x_address(4), B1 => lbl1_cx_n_8, B2 => x_address(4), ZN => lbl1_cx_n_10);
  lbl1_cx_count_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN298_lbl1_cx_n_7, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => x_address(2));
  lbl1_cx_g94 : MOAI22D0BWP7T port map(A1 => lbl1_cx_n_6, A2 => x_address(3), B1 => lbl1_cx_n_6, B2 => x_address(3), ZN => lbl1_cx_n_9);
  lbl1_cx_g95 : IND2D1BWP7T port map(A1 => lbl1_cx_n_6, B1 => x_address(3), ZN => lbl1_cx_n_8);
  lbl1_cx_count_reg_1 : DFKCNQD1BWP7T port map(CN => FE_PHN296_lbl1_cx_n_5, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => x_address(1));
  lbl1_cx_g97 : MOAI22D0BWP7T port map(A1 => lbl1_cx_n_4, A2 => x_address(2), B1 => lbl1_cx_n_4, B2 => x_address(2), ZN => lbl1_cx_n_7);
  lbl1_cx_g98 : IND2D1BWP7T port map(A1 => lbl1_cx_n_4, B1 => x_address(2), ZN => lbl1_cx_n_6);
  lbl1_cx_count_reg_0 : DFKCNQD1BWP7T port map(CN => FE_PHN283_lbl1_cx_n_3, CP => CTS_18, D => FE_DBTN23_memory_reset_out, Q => x_address(0));
  lbl1_cx_g100 : MOAI22D0BWP7T port map(A1 => lbl1_cx_n_2, A2 => x_address(1), B1 => lbl1_cx_n_2, B2 => x_address(1), ZN => lbl1_cx_n_5);
  lbl1_cx_g101 : IND2D1BWP7T port map(A1 => lbl1_cx_n_2, B1 => x_address(1), ZN => lbl1_cx_n_4);
  lbl1_cx_g102 : MOAI22D0BWP7T port map(A1 => lbl1_cx_n_1, A2 => x_address(0), B1 => lbl1_cx_n_1, B2 => x_address(0), ZN => lbl1_cx_n_3);
  lbl1_cx_g103 : IND2D1BWP7T port map(A1 => lbl1_cx_n_1, B1 => x_address(0), ZN => lbl1_cx_n_2);
  lbl1_cx_g104 : ND2D1BWP7T port map(A1 => x_increment_out, A2 => lbl1_cx_prev_incr, ZN => lbl1_cx_n_1);
  lbl1_cx_prev_incr_reg : DFD1BWP7T port map(CP => CTS_18, D => x_increment_out, Q => UNCONNECTED9, QN => lbl1_cx_prev_incr);
  lbl0_reg_n_layer_0_q_reg : EDFKCNQD1BWP7T port map(CN => FE_OFN5_FE_DBTN24_rst, CP => CTS_18, D => lbl0_n_500, E => lbl0_n_531, Q => lbl0_next_layer_0);

end routed;
