configuration counter5b_behaviour_cfg of counter5b is
   for behaviour
   end for;
end counter5b_behaviour_cfg;
