configuration reg_11_behaviour_cfg of reg_11 is
   for behaviour
   end for;
end reg_11_behaviour_cfg;
