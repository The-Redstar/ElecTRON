library IEEE;
use IEEE.std_logic_1164.ALL;

entity ge_register_tb is
end ge_register_tb;

