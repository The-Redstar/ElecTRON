configuration busy_counter_behaviour_cfg of busy_counter is
   for behaviour
   end for;
end busy_counter_behaviour_cfg;
